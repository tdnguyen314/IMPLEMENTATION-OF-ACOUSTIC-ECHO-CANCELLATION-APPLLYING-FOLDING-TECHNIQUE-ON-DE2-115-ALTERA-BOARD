--===========================================================--
--=================== Simulate the inputs ===================--
--===========================================================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;

entity Inputs_Simulation is
   port (
      RESET    : in  std_logic;
      SA_CLK   : in  std_logic;
      datax    : out byte_exdata;
      datad    : out byte_exdata);
end Inputs_Simulation;

architecture behavioural of Inputs_Simulation is
constant len : natural := 976;
type array_data is array(0 to len-1) of byte_data;
signal sdatax : array_data:=
--(others=>(others=>'0'));
("1111111111111111","0000000000000000","1111111111111111","1111111111111111","0000000000000000","0000000000000000","1111111111111111","1111111111111111","0000000000000000","1111111111111111","1111111111111111","0000000000000000","0000000000000000","1111111111111111","1111111111111111","0000000000000000","1111111111111111","1111111111111111","0000000000000001","1111111111111111","1111111111111110","0000000000000000","0000000000000001","1111111111111110","1111111111111111","0000000000000010","1111111111111110","1111111111111110","0000000000000010","0000000000000000","1111111111111101","0000000000000001","0000000000000001","1111111111111100","1111111111111111","0000000000000011","1111111111111101","1111111111111101","0000000000000100","0000000000000000","1111111111111011","0000000000000010","0000000000000011","1111111111111010","1111111111111111","0000000000000110","1111111111111100","1111111111111010","0000000000001000","0000000000000000","1111111111110101","0000000000000110","0000000000000111","1111111111110010","0000000000000000","0000000000001111","1111111111110010","1111111111110110","0000000000011011","1111111111110100","1111111111011110","0000000000111111","1111111111110110","1111111001110100","1111110111001000","1111111011110111","1111111110001110","1111111010001111","1111111011001110","0000000100101100","0000001010001110","0000000110101110","0000000010001001","1111111110101010","1111111001101010","1111111000100001","1111111110001110","0000000010000101","1111111111100110","1111111101111101","0000000001000011","0000000101100000","0000001001001011","0000001000111110","0000000001110110","1111111011000100","1111111101101101","0000000011011001","0000000010010110","1111111111001011","1111111111001100","1111111100011000","1111110110001110","1111110110011110","1111111101101010","0000000010011101","0000000010111010","0000000010010100","0000000000010111","1111111111011111","0000000010110111","0000000011101000","1111111100111001","1111111000110000","1111111100110000","1111111101110110","1111111001011100","1111111100000111","0000000101000011","0000000101010010","1111111110100000","1111111111011000","0000000110101000","0000001000001111","0000000100001010","0000000010001100","0000000011110110","0000000101110010","0000000100000110","1111111100100010","1111110100010010","1111110100000000","1111111010100110","1111111110101110","1111111101011011","1111111100011000","1111111111101010","0000000100010100","0000000100101111","0000000000100000","1111111101111110","0000000000101100","0000000011111000","0000000011011001","0000000001101011","1111111111111001","1111111100010000","1111111010001011","1111111101101011","0000000000100100","1111111100011010","1111111001000101","1111111110111111","0000000100110000","0000000000000011","1111111010101111","1111111111110010","0000000101010011","0000000001101100","1111111111000011","0000000011001110","0000000010010000","1111111010001110","1111111001011000","1111111111010110","1111111110100111","1111111010101100","1111111110111000","0000000011110100","1111111111110111","1111111100100100","0000000001010111","0000000011100100","1111111100100110","1111110110111011","1111111011000111","0000000011001100","0000000101001011","0000000000011111","1111111101110001","0000000001011110","0000000100010000","0000000001000111","1111111111100010","0000000011001011","0000000010101110","1111111100001110","1111111011011100","0000000001110110","0000000010110010","1111111100101111","1111111011010000","1111111111101011","0000000001001111","1111111110111011","1111111101101101","1111111101101101","1111111110110001","0000000010110111","0000000110001101","0000000011110111","0000000000100101","0000000001110100","0000000010100101","1111111110101011","1111111011000010","1111111010011111","1111111010101110","1111111101000100","0000000010011100","0000000100110110","0000000010001110","0000000001000011","0000000011001111","0000000011000100","1111111110111110","1111111011010001","1111111011010001","1111111110111111","0000000010111001","0000000011100101","0000000011001110","0000000011110001","0000000001101101","1111111110101011","0000000001101001","0000000100111100","1111111110000001","1111110110100010","1111111100100111","0000000101111011","0000000101100100","0000000101010001","0000001010011011","0000000111010001","1111111100001101","1111111011100010","0000000010100001","1111111110101001","1111110101110110","1111111001111110","0000000010100000","1111111110101100","1111111000101010","1111111111110101","0000001000110100","0000000011111100","1111111010101001","1111111010100010","1111111100110100","1111111001010110","1111111000100010","1111111110111111","0000000001100001","1111111100011011","1111111100000110","0000000011110111","0000000111001010","0000000001011110","1111111100100111","1111111101110111","0000000001100101","0000000100111010","0000000110010110","0000000011111001","0000000000001010","1111111111110000","0000000001010000","0000000001001001","0000000000001000","1111111111000010","1111111101101001","1111111110110101","0000000011011001","0000000101010001","0000000010010010","0000000000101000","0000000001001111","1111111110110110","1111111101000000","0000000010000010","0000000101101000","1111111110011111","1111110110100101","1111111001101111","0000000000110001","0000000001100001","1111111110111110","1111111101110101","1111111101100000","1111111110010101","1111111110111001","1111111100100010","1111111100101011","0000000011011101","0000000110011101","0000000000001010","1111111110000101","0000000101011000","0000000111110100","0000000011100111","0000000110110111","0000001110001000","0000001001111001","1111111111101010","1111111110001111","0000000001011101","0000000000000111","1111111110111110","0000000010011000","0000000101000010","0000000100111011","0000000101000100","0000000101101000","0000000110000000","0000000101110100","0000000010111010","1111111111110111","0000000010000000","0000000011111101","1111111110011010","1111111010001011","1111111111111100","0000000100101010","0000000000111000","0000000000000000","0000000011111111","1111111111101110","1111110111110111","1111111100001001","0000000011100100","1111111110100010","1111111001010011","0000000001001001","0000000111010110","0000000001000100","1111111100011101","0000000001001011","0000000100000010","0000000000110111","1111111110100111","1111111110011100","1111111101110001","1111111101110100","1111111110110111","1111111111000101","1111111101101011","1111111001110011","1111110110010011","1111111010000001","0000000011111110","0000001010010000","0000001000111001","0000000011101011","1111111101010001","1111111001000110","1111111010110000","1111111110110001","0000000000001101","1111111111110100","1111111110000101","1111111011011110","1111111100110001","0000000000110100","0000000000100011","0000000000110000","0000000111111101","0000001001110110","1111111110111000","1111111000110010","1111111111110000","0000000010000001","1111111011001100","1111111010111100","0000000000111000","0000000010000001","0000000010011101","0000000100101000","1111111111110101","1111111010011101","0000000001101100","0000001010000111","0000000101010010","1111111111010100","0000000010001110","0000000010101011","1111111110100010","0000000000110111","0000000101000000","0000000001010101","1111111110101111","0000000010101001","0000000001000011","1111111001101110","1111111011011011","0000000011011101","0000000010111100","1111111100111010","1111111101000111","0000000001001001","0000000010001110","0000000001011111","0000000000111011","0000000000110001","0000000001110011","0000000010000011","0000000000111011","0000000011101001","0000001000111111","0000001000001001","0000000011000000","0000000010001000","0000000000110000","1111111000101010","1111110100011101","1111111011010011","0000000000101101","1111111101000000","1111111010100111","1111111111001101","0000000010000000","1111111110001001","1111111001111100","1111111011100111","0000000001100101","0000000101100011","0000000011110001","1111111110011001","1111111001101000","1111111000100101","1111111100010011","0000000010000011","0000000101010110","0000000100111101","0000000001011000","1111111100000100","1111111011110111","0000000011011100","0000000110011010","1111111100110110","1111110100111111","1111111010100101","0000000010110010","0000000010100001","1111111110000111","1111111011111011","1111111110111000","0000000110101010","0000001001101100","0000000010101100","1111111110001111","0000000010101010","0000000011011100","1111111110001100","1111111101011111","1111111100110000","1111110110000000","1111110111100100","0000000100001000","0000000110010010","1111111101011111","0000000000011000","0000001011111010","0000001010110011","0000000001010010","1111111110110000","1111111111101010","1111111111001010","0000000010101000","0000000101110001","0000000001001101","1111111110110001","0000000110000010","0000001000110110","1111111110101010","1111110111011111","1111111110000010","0000000101001001","0000000010111111","0000000001001000","0000000101000010","0000000100100001","1111111100010000","1111111000001011","1111111100111101","0000000000001101","1111111100111010","1111111010101111","1111111101110100","0000000001000000","0000000000110101","1111111110111110","1111111100100100","1111111010000111","1111111010011100","1111111110110000","0000000010010100","0000000000010000","1111111011101010","1111111010011000","1111111010110100","1111111001101001","1111111011110101","0000000100000100","0000000111001000","1111111101011100","1111110101000010","1111111100100011","0000001001000100","0000000111011101","1111111100000011","1111111001100010","0000000000011010","0000000000111110","1111111010100011","1111111100010001","0000000101100111","0000000101010001","1111111011001101","1111111001111001","0000000011001001","0000000101111101","1111111110110111","1111111010010101","1111111100001110","1111111110000100","1111111101110010","1111111110001101","0000000000110011","0000000011100001","0000000001001111","1111111010001110","1111111000011001","1111111110011101","0000000000011110","1111111011001110","1111111010111110","0000000001001010","0000000011001000","0000000011001011","0000000111111111","0000000110111010","1111111001110100","1111110010100010","1111111011010011","0000000010101011","1111111100010111","1111110101000011","1111111001000000","0000000010011100","0000000110011010","0000000010111000","1111111111001010","0000000000110001","0000000001010100","1111111010100111","1111110110101000","1111111101011100","0000000011000011","1111111111010101","1111111110010111","0000000100011011","0000000100111010","1111111111110011","0000000000110001","0000000011000110","1111111100101110","1111110110011111","1111111001111110","1111111110110101","1111111110010111","1111111110100110","0000000001100110","0000000010000110","0000000000001101","0000000001000111","0000000110100001","0000001100100000","0000001100011000","0000000100100111","1111111101101100","1111111110101001","0000000010011000","0000000001110011","1111111111000111","1111111111001101","0000000001111001","0000000011111100","0000000010110111","1111111110010111","1111111001010101","1111110111100111","1111111011010110","0000000010001101","0000000100101010","1111111111001011","1111111010000000","1111111100001101","1111111111001011","1111111110011001","0000000001111100","0000001010010100","0000001010101101","0000000010101100","0000000000000011","0000000011010011","0000000001101011","1111111101010101","1111111101110101","1111111110101101","1111111100101100","1111111110100001","0000000011001011","0000000001100110","1111111101100011","0000000000001110","0000000011100000","1111111111011001","1111111010000001","1111110111001011","1111110010111000","1111110011110111","0000000000100110","0000001001010100","0000000010000100","1111111011101011","0000000001101110","0000000101010010","0000000000101010","0000000000110100","0000000011001111","1111111100011100","1111110110101100","1111111101101001","0000000100011111","0000000000101110","1111111100011011","1111111101101101","1111111111010101","0000000000101001","0000000010011010","0000000000111101","1111111110001101","1111111111001011","0000000001000011","0000000000000101","1111111101110101","1111111011001000","1111111001010010","1111111010100100","1111111011010001","1111111011001011","0000000011110110","0000010000110111","0000001101011111","1111111011100010","1111110100000111","1111111011000101","1111111111111011","0000000000100000","0000000001100001","1111111101111101","1111111001010001","1111111110001010","0000000100101110","0000000000101111","1111111011011101","1111111101110111","1111111111101101","1111111110110110","0000000001110110","0000000011000011","1111111101010100","1111111011110100","0000000001111011","0000000001111001","1111111010010111","1111111001000011","1111111110010011","1111111111111100","1111111111001110","0000000001010001","0000000001101100","1111111110011110","1111111110111010","0000000011111101","0000000011111100","1111111100111011","1111111001111111","1111111110111100","0000000000111111","1111111101110010","0000000010010100","0000001101110111","0000001101000101","1111111110011001","1111110110110101","1111111011011111","1111111110000101","1111111101001101","0000000000010101","0000000001111110","1111111101110111","1111111100101101","1111111111001111","1111111100100011","1111111001100011","0000000000011001","0000001000100111","0000000110010001","0000000001100011","0000000101111111","0000001011111100","0000000111010100","1111111110100000","1111111111001101","0000000101110011","0000000100101100","1111111110000100","1111111110001110","0000000010011110","0000000000110111","1111111101101011","1111111110101011","1111111100011010","1111110100111001","1111110011010100","1111111010000011","0000000000001000","0000000010101101","0000000011011011","0000000000010100","1111111010001011","1111110110000001","1111110111001100","1111111110111101","0000001000011011","0000001001001010","0000000010000101","1111111111011001","0000000001101001","0000000000000010","1111111101000000","1111111110010011","1111111111111011","1111111111011101","1111111110110110","1111111100001101","1111111010100010","0000000000010100","0000000110000011","0000000011010100","0000000001011100","0000000100001010","0000000000111110","1111111101011101","0000000101101010","0000001011100011","0000000011000001","1111111101101001","0000000010101111","0000000001101110","1111111100001101","1111111111010111","0000000001100011","1111111100010101","1111111110011100","0000000100100000","1111111101001010","1111110100101100","1111111100010110","0000000011100011","1111111110111000","1111111111101100","0000000111010011","0000000011011111","1111111010001011","1111111011010000","1111111110000111","1111111010000101","1111111001111110","0000000000001011","0000000010010011","0000000000110001","0000000000011011","1111111110110010","1111111101110101","0000000001001111","0000000010010100","1111111111010011","0000000001011001","0000000101101010","0000000000011010","1111111000011000","1111111010100110","0000000001100001","0000000100100010","0000000101111100","0000000011010110","1111111001010111","1111110101000011","1111111111000000","0000000110001110","1111111110010111","1111110110111011","1111111100111010","0000000100110101","0000000010011000","1111111010110000","1111110111110011","1111111011011000","0000000000111101","0000000011000011","0000000000101001","1111111110010101","0000000000001111","0000000100001100","0000000011011110","1111111011111111","1111110110010100","1111111010100110","0000000001110110","0000000001100011","1111111110101000","0000000001000011","0000000010111111","0000000000100000","0000000001000110","0000000011110010","0000000000000101","1111111101010101","0000000101101001","0000001011111110","0000000011011011","1111111010100010","1111111111011101","0000000110100001","0000000011100000","1111111101110000","1111111101001100","1111111110001110","1111111110000000","1111111111100100","0000000011011111","0000000101011110","0000000010101110","1111111101111001","1111111011010110","1111111011000000","1111111010000101","1111111001001111","1111111010111100","1111111110110011","0000000010010111","0000000100000000","0000000100001101","0000000101011101","0000000111011111","0000000101101011","0000000000011110","1111111110010000","1111111101111000","1111111001111110","1111111000110000","0000000000011100","0000000110001001","0000000001100110","1111111110000011","0000000001111010","0000000010101011","1111111110001000","1111111101110110","0000000000011100","1111111111001100","1111111110111101","0000000011000011","0000000011101110","0000000000001011","0000000001001110","0000000110100010","0000000111100100","0000000010110001","1111111110001011","1111111110101010","0000000010010110","0000000001011111","1111111011111001","1111111100011101","0000000010100010","1111111111000100","1111110101001010","1111111000011100","0000000100001011","0000000011101001","1111111100011001","1111111110011010","0000000001000110","1111111100000100","1111111100010110","0000000011101011","0000000010011101","1111111011111101","1111111110001011","0000000001010100","1111111100011001","1111111100001000","0000000100110001","0000000101111110","1111111101010010","1111111010010110","1111111111100011","0000000010100011","0000000001100100","0000000000101110","0000000000010111","0000000000010001","0000000001011001","0000000011100001","0000000101100000","0000000100000101","1111111110001000","1111111011011100","0000000001100100","0000000111010010","0000000100010101","0000000000110010","0000000100101101","0000001001011011","0000000111100011","0000000010111101","0000000001111011","0000000010110101","1111111111001000","1111110111000111","1111110110000100","0000000000000001","0000000100010100","1111110111111101","1111101110001111","1111111001110111","0000001001011110","0000000101001101","1111111000001010","1111111001110100","0000000100011110","0000000100010010","1111111100000011","1111111100100011","0000000101000101","0000000110110110","1111111110110111","1111111000000111","1111111001000111","1111111101011100","1111111110000101","1111111010011101","1111111001111101","0000000001100000","0000001001011111","0000001000100111","0000000010011111","1111111110111101","1111111101100111","1111111100111111","1111111111001101","0000000010010111","0000000011001111","0000000011011000","0000000001100001","1111111011000011","1111110111011110","1111111101101010","0000000100110100","0000000100010110","0000000001110001","0000000001010011","0000000000001010","0000000000000010","0000000001011010","1111111110010101","1111111001110000","1111111101010001","0000000100010001","0000000100101000","0000000001100011","1111111111100001");
--("0000000000000000","0000000000000000","1111111111111111","1111111111111111","0000000000000000","1111111111111111","0000000000000000","1111111111111111","1111111111111111","0000000000000000","1111111111111111","1111111111111111","0000000000000000","0000000000000000","1111111111111111","1111111111111111","0000000000000000","1111111111111111","1111111111111111","0000000000000000","0000000000000000","1111111111111111","1111111111111111","0000000000000000","1111111111111111","1111111111111111","0000000000000000","0000000000000000","1111111111111111","0000000000000000","0000000000000000","1111111111111111","1111111111111111","0000000000000000","0000000000000000","1111111111111110","0000000000000000","0000000000000001","1111111111111110","1111111111111111","0000000000000001","1111111111111111","1111111111111110","0000000000000010","0000000000000000","1111111111111100","0000000000000000","0000000000000011","1111111111111100","1111111111111101","0000000000000101","1111111111111111","1111111111111010","0000000000000100","0000000000000011","1111111111111000","0000000000000000","0000000000001000","1111111111111001","1111111111111010","0000000000001100","1111111111111111","1111111111101011","0000000000100011","0000000011100011","0000001000000001","0000001001010010","0000000011000011","1111111011010111","1111111100101101","0000000011010100","0000000011010100","1111111110101010","1111111101101011","1111111100000100","1111110110111001","1111111000110111","0000000010001011","0000000010101000","1111111010001011","1111111001001001","1111111110101100","1111111110110110","1111111110100110","0000000101100000","0000001010011100","0000000111101111","0000000101011111","0000000101000100","0000000000101010","1111111100100100","1111111111010001","0000000011111100","0000000100100011","0000000010101001","0000000001000101","0000000001011000","0000000011110010","0000000100111100","0000000010011111","0000000000001100","0000000001010001","0000000011001111","0000000010101100","1111111111001000","1111111100000001","1111111110010101","0000000011111010","0000000100001111","1111111111110010","0000000000000011","0000000101111011","0000001001001100","0000001000000100","0000000111100000","0000001000011101","0000000110111010","0000000000010111","1111111001111000","1111111011101000","0000000001101011","0000000000000100","1111111010110111","1111111111010011","0000000110001111","0000000001110110","1111111100010001","0000000000111110","0000000011010101","1111111100111001","1111111100110110","0000000100001111","0000000010101001","1111111010111011","1111111100101111","0000000100011011","0000000101101011","0000000001111111","1111111111011101","1111111111100010","0000000010011010","0000000100011001","0000000001101010","1111111111101100","0000000010010011","0000000010010111","1111111110011000","1111111110011010","0000000001011101","0000000000110000","1111111111010111","1111111111111111","1111111101110101","1111111011111001","0000000001011001","0000000111011111","0000000101010111","0000000001001111","0000000001001111","0000000001111110","0000000011100101","0000000101110011","0000000000011011","1111110111000001","1111111001111000","0000000100000101","0000000000111001","1111110110110000","1111111011100000","0000000110101000","0000000011111001","1111111101100100","0000000010111000","0000000110000101","1111111101010011","1111111010101001","0000000100011011","0000000110001110","1111111011110000","1111111001010011","0000000010000011","0000000100101001","1111111110101001","1111111100100011","0000000000000010","0000000010110110","0000000101101000","0000001001000000","0000000111011011","0000000000100100","1111111100010101","1111111101011000","1111111110001110","1111111110000001","0000000001010101","0000000100110110","0000000001010110","1111111101001100","0000000010101001","0000000111111111","1111111111110110","1111110111100001","1111111111001101","0000000111001000","1111111101111100","1111110100010001","1111111011100100","0000000110001011","0000000110011001","0000000100010100","0000000101000010","0000000011001101","0000000001001100","0000000011110011","0000000101110101","0000000011011100","0000000001000000","0000000001010001","0000000011101110","0000000111100010","0000001000100010","0000000100010010","1111111111101001","1111111101001101","1111111010011101","1111111010011010","0000000000101010","0000000101110111","0000000011100000","0000000000110101","0000000101010100","0000001010101101","0000001000001101","0000000001100101","0000000000110101","0000000100000001","1111111111001111","1111110100111111","1111110101101001","1111111110111110","1111111110101011","1111111000110001","1111111110010111","0000000101111111","1111111111101001","1111111000111100","1111111110100000","0000000001101110","1111111110010100","0000000011011101","0000001011010110","0000000100111010","1111111010011111","1111111010100110","1111111010111001","1111110111000010","1111111100001010","0000000101100010","0000000010111110","1111111100100100","0000000001001001","0000001001010000","0000001011000110","0000001001001110","0000000010111011","1111111001001011","1111111000001010","0000000000100110","0000000010111000","1111111110010000","1111111111101001","0000000100000010","0000000010011000","0000000001110000","0000000110010011","0000000100111110","1111111100111100","1111111010111100","1111111110101110","1111111110100110","1111111100010000","1111111100011111","1111111101000011","1111111111000111","0000000011110001","0000000010100001","1111111010001000","1111111000001011","1111111111011000","0000000010111010","0000000000010000","1111111110010011","1111111011101001","1111111001010000","1111111111000001","0000000110011000","0000000001000000","1111110110100001","1111110111001111","1111111110011011","0000000001100111","0000000100000001","0000000110010000","0000000010010101","1111111101010101","1111111110110000","0000000000101000","1111111110101110","1111111111010000","0000000001110110","0000000000000001","1111111100101101","1111111100101100","1111111100011000","1111111010101001","1111111011010010","1111111101101000","0000000000111011","0000000110101100","0000001000101101","0000000001101111","1111111100001101","1111111111001111","1111111111100111","1111111001010111","1111111010010100","0000000011100001","0000000100110011","1111111100011110","1111110111100000","1111111001010000","1111111110001011","0000000100101010","0000000101001011","1111111100000110","1111110111001000","1111111101010010","1111111111010000","1111111000000110","1111110111101000","1111111101110011","1111111010110010","1111110011110011","1111110111010001","1111111100100101","1111111001110000","1111111010000101","0000000001011010","0000000010100110","1111111110110001","0000000010010100","0000000111111101","0000000101011111","0000000001010101","0000000001110001","0000000010010111","0000000011001110","0000000110001100","0000000100010100","1111111100110011","1111111010000110","1111111101001101","1111111101100110","1111111011110110","1111111100010010","1111111100010011","1111111101000010","0000000011101011","0000001001110011","0000000101110101","1111111111000101","0000000001011100","0000000111110010","0000000111000100","0000000010010001","0000000010001110","0000000100111011","0000000011110000","0000000000100111","0000000000100111","0000000001101010","0000000000011000","1111111111000001","1111111110110011","1111111110010000","0000000001010110","0000001010111010","0000010000001110","0000000111101010","1111111011111010","1111111100000111","0000000011110100","0000000100000100","1111111010100110","1111110011101010","1111111000010101","0000000001111010","0000000100001100","0000000000010000","1111111110101001","1111111110000010","1111111011100011","1111111110101001","0000000111001101","0000000110111001","1111111100110111","1111111001110111","0000000010010010","0000001010011111","0000001011110010","0000000110010011","1111111101111110","1111111100010111","0000000001110101","0000000001011000","1111111011101111","1111111111000101","0000000110001000","0000000001101000","1111111001100110","1111111011110010","0000000001010101","0000000010111111","0000000101001010","0000000101111111","0000000010001011","0000000000010010","0000000000001111","1111111100001000","1111111011101110","0000000011001111","0000000011011101","1111111011000011","1111111110010001","0000001010001101","0000000111001110","1111111001011001","1111110111001101","1111111110110011","0000000001100110","0000000000110110","0000000001010000","1111111110100011","1111111000111111","1111111000101011","1111111111101111","0000000101010001","0000000001100010","1111111011110111","0000000000010101","0000000111001100","0000000000001110","1111110100001100","1111110101110100","1111111110001101","1111111111111101","0000000001011111","0000000100111101","1111111111011011","1111110110111001","1111111010011001","0000000011001111","0000000110001010","0000000110111110","0000000101000011","1111111100101000","1111111001010011","1111111111110000","0000000000001000","1111111000110100","1111111001010010","1111111110101011","1111111110101001","0000000000101010","0000000110100010","0000000011101101","1111111100110110","0000000000010110","0000000110101111","0000000100110010","0000000001000100","1111111110111100","1111111010100001","1111111001111110","0000000000010111","0000000010111011","1111111111011101","1111111110011001","1111111110110101","1111111101110010","1111111111101101","0000000010010101","0000000000110101","0000000001111101","0000000111010110","0000000101100001","1111111100111000","1111111001100100","1111111011001000","1111111100010000","0000000000000100","0000000011110011","0000000000100010","1111111100011001","1111111100101000","1111111000101110","1111110010001101","1111110111100011","0000000100101110","0000000111000111","1111111110010011","1111111000011011","1111111010000010","1111111110011101","0000000001101010","0000000001111101","0000000010000100","0000000100101011","0000000100010110","1111111101001001","1111110111100101","1111111010100100","1111111110110011","1111111101111100","1111111110101101","0000000101110110","0000001010000101","0000000100000011","1111111101011101","0000000001000000","0000000110100110","0000000011011000","1111111111001100","0000000011101010","0000001001000010","0000000111110100","0000000100111101","0000000001010001","1111111011011011","1111111101110001","0000001000011110","0000000110010000","1111110110101101","1111110110111000","0000000111011111","0000001000000011","1111111000001011","1111110111101010","0000000101100000","0000000110010000","1111111100011000","1111111100001000","0000000001011001","0000000000001011","1111111101101001","1111111110001001","1111111101000011","1111111100100010","1111111111000010","1111111110011000","1111111100110001","0000000011100110","0000001011010111","0000000111000101","1111111110111010","1111111111110010","0000000101001110","0000001000000100","0000000111100110","0000000001010000","1111111001011001","1111111011101010","0000000010001100","1111111110100001","1111111001110110","0000000000001100","0000000010111100","1111111010010101","1111111001001111","0000000010010000","0000000010011100","1111111101101001","0000000010001110","0000000100001100","1111111010111000","1111111000011111","0000000000100000","1111111111001001","1111110110011001","1111111000100010","0000000001001011","0000000011101110","0000000011011000","0000000010011001","1111111110010100","1111111110111011","0000000101001100","0000000010011001","1111111000101111","1111111100001100","0000001000110000","0000001001001001","0000000001000101","0000000001011011","0000000101000000","1111111111110110","1111111000000100","1111110110000001","1111110111000111","1111111010101101","0000000001011111","0000000011110000","1111111110111010","1111111110100010","0000000101111000","0000000111101010","0000000000100111","1111111101100100","0000000001010011","0000000011101010","0000000111000010","0000001101111100","0000001010111101","1111111011010111","1111110110001001","0000000010000010","0000000101001001","1111110111100000","1111110011110010","0000000001110111","0000000111111100","1111111101111100","1111111001101111","0000000001100101","0000000011111000","1111111101010110","1111111100100110","0000000010110000","0000000100000101","0000000001010100","0000000011001010","0000000110011101","0000000100000110","1111111111100101","1111111101010010","1111111011011011","1111111100010001","0000000010001100","0000000100101111","0000000000010101","0000000000010101","0000000110011010","0000000100010001","1111111010101111","1111111001100000","1111111111011000","0000000001000100","0000000001010111","0000000011001000","1111111111110010","1111111100111100","0000000100011110","0000001001100010","0000000000000100","1111111000010010","1111111101010011","1111111111010011","1111111001011010","1111111011110011","0000000100011010","0000000001100000","1111111000010110","1111111010011011","0000000010100011","0000000010010111","1111111110000110","1111111111101100","0000000010110110","0000000001000100","1111111110111110","0000000010001100","0000000111001111","0000001000100011","0000000101111011","0000000010001100","0000000000001111","0000000001101111","0000000100011111","0000000101010010","0000000101001111","0000000101100010","0000000011111000","0000000010100000","0000000110000111","0000001000100010","0000000010001010","1111111011110011","1111111110000000","1111111111010110","1111111011000110","1111111100110110","0000000100001100","0000000010001101","1111111000010111","1111110101001101","1111111010000001","0000000000000000","0000000011111010","0000000001001001","1111111001111101","1111111100010100","0000000111000111","0000001000000110","0000000001010010","0000000100111011","0000001101001100","0000001000101110","1111111110110100","1111111100111010","1111111100001010","1111110111101110","1111111000100001","1111111101111000","1111111101110010","1111111010111100","1111111100101110","1111111111011101","1111111111110011","0000000000110001","1111111111000101","1111110110101100","1111110010011001","1111111100111011","0000001010101000","0000001010011101","0000000010010000","0000000001111100","0000000110010101","0000000010001001","1111111001100011","1111111011101110","0000000111011001","0000001100100011","0000000101000101","1111111010111101","1111111000011001","1111111100010011","1111111110110110","1111111101001000","1111111100101100","0000000001001100","0000000101011010","0000000100010100","0000000001010111","0000000000100011","0000000000001110","1111111111011110","0000000000011110","0000000010101110","0000000011101111","0000000100001000","0000000100110011","0000000010110110","1111111100100000","1111110110101111","1111111000001111","1111111111100101","0000000100001111","0000000010011000","1111111110111011","1111111110101110","0000000000100011","0000000001100010","0000000000100010","1111111110000000","1111111100111001","1111111111101010","0000000010100010","0000000000111101","1111111110011110","0000000000101011","0000000100011110","0000000011110000","0000000000000100","1111111110110110","0000000001001010","0000000100101100","0000000111011111","0000000111000001","0000000001001100","1111111001100011","1111111000010000","1111111110011010","0000000010001000","1111111110111110","1111111110101101","0000000101010100","0000000110101110","1111111111101000","1111111111000100","0000000110110110","0000000100101111","1111111001000111","1111111010001011","0000000111000110","0000001000001101","1111111101101111","1111111100001000","0000000001010100","1111111110111110","1111111100101010","0000000100011001","0000001001010001","0000000011100011","0000000001001000","0000000101100011","0000000011110011","1111111110100000","0000000010110000","0000001001111010","0000000111000010","1111111111110110","1111111100110010","1111111011100001","1111111101010101","0000000100010011","0000000110011110","1111111110011000","1111110111111000","1111111010010011","1111111110110100","0000000001010111","0000000010110100","0000000001011010","1111111111001000","1111111111110001","1111111111110101","1111111111000000","0000000011100001","0000001000001001","0000000100001110","0000000001001101","0000000110100110","0000000111000011","1111111111110000","0000000001001000","0000001000011000","0000000101000010","1111111111100010","0000000100000000","0000000011110101","1111111001011100","1111111001110100","0000000110001010","0000000111000100","1111111101000011","1111111011011110","1111111111111001","1111111110111000","1111111101110011","0000000000001101","1111111110000110","1111111001010010","1111111011010111","0000000000110011","0000000000011100","1111111100001001","1111111010010100","1111111011111001","1111111111010110","0000000011000010","0000000100001011","0000000010000111","1111111111101100","1111111110111100","1111111110100111","1111111110000011","1111111111110001","0000000011110101","0000000100000011","1111111110000100","1111111010001110","1111111101101001","0000000000111110","1111111111001101","1111111110000101","1111111111101000","1111111110101100","1111111011101011","1111111011010100","1111111101011011","0000000010000100","0000001010100000","0000001111010001","0000001000011011","1111111110010111","1111111101010110","0000000000110101","1111111111000010","1111111011001000","1111111011101101","1111111110010000","1111111111001101","1111111111101001","1111111111001100","1111111101010110","1111111110000111","0000000001011001","1111111110111101","1111110110011000","1111110100110010","1111111110111001","0000000110011000","0000000010000101","1111111100111100","1111111111110111","0000000010110110","0000000000111111","0000000010001100","0000000110001101","0000000001100111","1111110111001101","1111110110100011","1111111110100100","0000000000000010","1111111010010001","1111111001000101","1111111101011110","1111111111111000","1111111111001111","1111111110111011","1111111111110110","0000000001000101","0000000000110011","1111111111011000","0000000000011101","0000000001110010","1111111100001101","1111110101000111","1111111000101000","0000000001000001","0000000000101101","1111111011101000","1111111010111101","1111111100101011","0000000000110101","0000001000100110","0000001000010001","1111111101010110","1111111100000101","0000000111011110","0000001000001110","1111111101110010","1111111101101100","0000000011011101","1111111110110011","1111111010111100","0000000010110011","0000000111100110","0000000011010001","0000000001111011","0000000011000010","0000000000000110","1111111111101101","0000000001110001","1111111100110101","1111110111111010","1111111100111111","0000000001011110","1111111111000110","0000000000100100","0000000100100000","0000000001001100","1111111111001111","0000000101101000","0000000110101001","1111111110110011","1111111101011001","0000000011110010","0000000110110010","0000000110010011","0000000100110010","0000000000111101","0000000001111011","0000001001001111","0000000111011101","1111111011101101","1111111001101110","0000000000101000","1111111110110001","1111111011110010","0000000101110011","0000001011101011","1111111110101100","1111110100101011","1111111110000111","0000000111100000","0000000001010010","1111111001010110","1111111011111110","0000000000100011","1111111110010111","1111111010101111","1111111100110110","0000000001010101","0000000000111010","1111111101110100","0000000000001011","0000000110011001","0000000110111111","0000000001111001","1111111111110011","0000000001011110","1111111111110010","1111111011001100","1111111011101000","0000000001001101","0000000010011110","1111111101010011","1111111011100101","0000000000011100","0000000000111010","1111111001110001","1111111000000101","0000000000110101","0000000111101110","0000000110010110","0000000011101101","0000000010110111","0000000001001100","0000000000010000","0000000001010100","0000000001111011","0000000011001011","0000000101110011","0000000100101011","1111111111011111","1111111100101111","1111111100111000","1111111100011001","1111111101100011","0000000000011010","0000000000001100","1111111111001100","0000000001010000","1111111111111100","1111111010010110","1111111100010100","0000000101000100","0000000101010001","1111111101010110","1111111011000100","1111111111010011","0000000100010101","0000001010011011","0000001100100110","0000000101110101","0000000001011010","0000000110100101","0000000111111011","0000000000111001","1111111111111010","0000000100110100","0000000010100101","1111111110110110","0000000011110001","0000000111011100","0000000011100111","0000000010011000","0000000100100100","0000000010111110","0000000001100001","0000000000110010","1111111010000001","1111110111000011","0000000001010101","0000000101111001","1111111010100011","1111110110110001","0000000000110001","0000000000010101","1111110111001001","1111111011011010","0000000011101101","1111111111011001","1111111101011001","0000000101000101","0000000011101111","1111111010110000","1111111011111101","1111111111001011","1111111001101001","1111111011000110","0000000110110011","0000000111111001","1111111110110001","1111111101111111","0000000010110100","0000000010100111","0000000000111000","1111111101010100","1111110101011001","1111110101100011","0000000000110110","0000000100100100","1111111101111000","1111111101010100","0000000000101110","1111111101110111","1111111110001101","0000000100110001","0000000010010011","1111111010010111","1111111101110111","0000000011101010","1111111101111100","1111111010101100","0000000001101111","0000000001110001","1111111000110001","1111111000010100","1111111111101000","0000000011000010","0000000101100100","0000001000100000","0000000011010001","1111111001000100","1111110100010010","1111110101111011","1111111111000100","0000001101010110","0000001101101101","1111111011000001","1111110010001010","0000000000011001","0000001010110001","0000000010101111","1111111011010000","1111111101111100","0000000000110010","0000000000110001","0000000000000110","1111111101010001","1111111011101110","1111111101101000","1111111100101110","1111111010100100","1111111111100010","0000000101110000","0000000100011010","0000000010011010","0000000011110111","0000000001001110","1111111101010011","0000000000100010","0000000011010101","1111111110001110","1111111010010010","1111111011010111","1111111001111000","1111111001100001","0000000010001101","0000001001001000","0000000001111101","1111110111100010","1111111000110010","1111111111011100","1111111110010010","1111111000100010","1111111010010001","0000000010111000","0000000110110011","0000000011101110","0000000010010100","0000000100110001","0000000101001001","0000000010110101","0000000000111111","1111111110000011","1111111010000000","1111111010110001","0000000001000000","0000000101100000","0000000100011001","0000000000001011","1111111100011010","1111111011110101","1111111110110000","0000000001111010","0000000010101010","0000000010000000","0000000010001101","0000000100000100","0000000100101010","1111111111101100","1111111001110010","1111111110000011","0000001001101010","0000001100001011","0000000011001011","1111111101011010","1111111111100101","0000000000101000","1111111111101110","0000000001110111","0000000010001010","1111111100111100","1111111010110111","1111111111010101","0000000001011100","1111111111110101","0000000001100000","0000000011110111","0000000010000100","0000000010101111","0000000111111000","0000000111011011","0000000010001110","0000000011111111","0000001001000011","0000000110001110","0000000000101100","1111111111101001","1111111101010100","1111111010001010","1111111110001110","0000000011001111","0000000000011100","1111111110111011","0000000100000010","0000000011111100","1111111101011111","1111111101101111","0000000011001010","0000000001111111","1111111100000001","1111111000111110","1111111000100111","1111111001100111","1111111011011111","1111111011100001","1111111011011000","1111111110000100","0000000000001001","0000000001100000","0000000111001010","0000001010001000","0000000000100011","1111110110000010","1111111001110000","0000000010001011","0000000000110011","1111111011111010","1111111110101111","0000000101101101","0000000111001001","0000000001011010","1111111100100111","1111111111000011","0000000001100101","1111111101001001","1111111011111110","0000000100111110","0000001001101000","0000000011100001","0000000001101110","0000000101011000","1111111111110011","1111111000101001","1111111111100100","0000000110000010","1111111101001111","1111111000101100","0000000101001010","0000001100001111","0000000010111100","1111111101110101","0000000011000111","0000000000100001","1111110110001100","1111110111101001","0000000011001011","0000000100111010","1111111100010011","1111111001101011","1111111111000010","0000000001101000","0000000000110000","0000000001001110","1111111111011100","1111111010000101","1111111001110010","1111111111011000","1111111111110111","1111111010001000","1111111000101100","1111111101011101","0000000001101100","0000000011101011","0000000100001001","0000000010101000","0000000010001000","0000000011101101","0000000010011001","1111111111010001","0000000000011111","0000000010000110","1111111110011010","1111111100110000","0000000001100011","0000000011100000","0000000000010000","1111111111111111","0000000000101001","1111111100011010","1111111010100001","1111111110110110","1111111111110010","1111111101101111","0000000011110011","0000001100001111","0000000111110100","1111111011001001","1111110110001001","1111111011111010","0000000100100110","0000000111011000","0000000000001101","1111111000001100","1111111011100011","0000000100010001","0000000101001101","0000000010011000","0000000011011110","0000000001110100","1111111011110011","1111111110000111","0000001000011001","0000001001011100","1111111111111001","1111111101000101","0000000100100010","0000000111100101","0000000001001111","1111111011111011","1111111100001001","1111111100010011","1111111100111011","0000000011000111","0000001000110111","0000000101101100","0000000000010001","0000000000100011","1111111111110011","1111111100000110","0000000000100111","0000001010001100","0000000111100011","1111111100011000","1111111011001100","0000000001111011","0000000010110100","1111111111010111","1111111101101000","1111111010111001","1111111000000101","1111111010000010","1111111110001010","0000000000101000","0000000010000000","0000000000110111","1111111110000010","1111111110110111","0000000000111010","1111111111011111","0000000001010001","0000000111110010","0000000110000011","1111111101101100","0000000000101011","0000001010011110","0000000101111000","1111110111100011","1111110100000010","1111111010011111","1111111110010011","1111111110000001","1111111100100100","1111111100110011","0000000011000101","0000001000100100","0000000001101001","1111111000100101","1111111110101010","0000001000101110","0000000100010110","1111111100011100","0000000000000101","0000000100101010","0000000000011100","1111111101110000","0000000001110000","0000000101110110","0000001001110001","0000001100101101","0000000110010010","1111111011110111","1111111100011011","0000000010100110","0000000001011101","0000000000010111","0000000100110001","0000000010100011","1111111011101111","1111111111011010","0000000100011000","1111111101001011","1111111010100000","0000000101001011","0000000110011110","1111111011010001","1111111011001011","0000000010001010","1111111110000110","1111111100111000","0000001000101010","0000001010000110","1111111101100111","1111111101101000","0000000110110011","0000000010011000","1111111011100001","0000000001110111","0000000011110000","1111111001110101","1111111001000110","0000000010011110","0000000010110110","1111111110011001","0000000010010101","0000000110000111","0000000010000110","1111111111110101","0000000010010000","0000000010000101","0000000000100001","0000000001110100","0000000010010100","1111111111110100","1111111101110111","1111111101110110","1111111111000110","0000000000111011","1111111111111010","1111111010101101","1111110111010000","1111111010011010","1111111111110100","0000000001000000","1111111111010011","0000000000111000","0000000101011111","0000000101100000","0000000000011000","1111111111100001","0000000011100000","0000000000110110","1111110111111000","1111110111100100","0000000010000111","0000001001000100","0000000111110100","0000000110101101","0000000110010001","0000000001001000","1111111100001010","1111111110100100","0000000010010011","1111111111110100","1111111110001001","0000000100110100","0000001010001110","0000000011101100","1111111010110011","1111111101010101","0000000101001110","0000000101100000","0000000000101100","1111111111010001","1111111111110000","1111111110010111","1111111101000010","1111111101011010","0000000000000001","0000000110000001","0000001010010111","0000000110001100","0000000000001101","0000000100000011","0000001100010001","0000001011011110","0000000011111111","0000000001011001","0000000101101001","0000001001110011","0000000111011110","1111111110101001","1111111001000010","1111111110010000","0000000100100110","0000000000010011","1111111001010011","1111111010011111","1111111101001010","1111111011100101","1111111110010011","0000000110110111","0000001010011010","0000000110110010","0000000010110001","1111111111110000","1111111110100110","0000000010001100","0000000101011101","0000000011001001","0000000001101001","0000000011101111","0000000000010010","1111111000000000","1111111000100101","0000000010011011","0000000111001100","0000000011101001","0000000010000010","0000000110000010","0000001000111111","0000000111010011","0000000101000001","0000000100101100","0000000010101100","1111111111000010","0000000000101011","0000000110110010","0000000110110000","0000000001000000","0000000000110011","0000000100111011","0000000010111010","1111111101000011","1111111011111101","1111111111000001","0000000011001000","0000000110001111","0000000010101100","1111111010111100","1111111010110110","0000000000110111","0000000001001010","1111111111110010","0000000100100011","0000000101001000","1111111100100010","1111111001110000","0000000000010000","0000000001110110","1111111110100001","0000000000001100","0000000010001001","1111111111110010","0000000001100010","0000000101001111","1111111110101010","1111110101011101","1111111010000000","0000000011100000","1111111111111111","1111110101110100","1111110110000111","1111111111101101","0000000101010011","0000000010110111","1111111110110011","1111111100010011","1111110111100111","1111110010010000","1111110110000000","0000000001100000","0000000100110100","1111111101110000","1111111011111111","1111111111100110","1111111001110000","1111110001101110","1111111011001000","0000001011010011","0000001000101000","1111111001000001","1111110101011001","1111111111100110","0000000110111001","0000000100101010","1111111111000101","1111111100110001","1111111110011111","0000000001000000","0000000100100000","0000001010011010","0000001001000110","1111111000111100","1111101100100100","1111111000010101","0000001010010010","0000000110110100","1111111001010101","1111111010000110","0000000001101100","0000000001000011","1111111111110101","0000000011010100","0000000001000110","1111111011010111","0000000000000110","0000001001001001","0000000101010101","1111111010100011","1111111011000101","0000000100001110","0000000100110100","1111111100001011","1111111010000110","0000000010101110","0000000111011010","0000000000100101","1111111010000001","1111111011101100","1111111101100000","1111111100010101","1111111111000110","0000000010001111","1111111101110000","1111111001111001","1111111110100001","0000000001011001","1111111110101101","0000000010000100","0000001001010111","0000000111100101","0000000010011001","0000000100001000","0000000100000001","1111111101101010","1111111101001010","0000000010101101","0000000011011011","0000000011000000","0000000101110100","0000000001111001","1111111000110001","1111111010001010","0000000010111001","0000000100010100","0000000010010010","0000000100100110","0000000100101111","0000000001100110","0000000010110011","0000000100001011","1111111111001001","1111111011100101","1111111110011000","1111111111101001","1111111101101100","1111111110011100","0000000000000110","1111111101110111","1111111010001111","1111111001110000","1111111110000101","0000000100100101","0000000101011010","1111111111000010","1111111100000101","0000000000011010","0000000001100100","1111111100010100","1111111001100001","1111111011011110","1111111110000001","0000000000100101","0000000001010000","1111111101111100","1111111100001110","1111111101111111","1111111100100001","1111111011010000","0000000010011010","0000000111010000","1111111111010001","1111111001111110","0000000001010101","0000000011101110","1111111100000111","1111111101101100","0000000110100100","0000000011011011","1111111100010100","0000000001001101","0000000100100010","1111111100111000","1111111100000100","0000000010111011","1111111100110101","1111110010010010","1111111001111111","0000000110001001","0000000001100000","1111111010111000","0000000001000010","0000000101000111","1111111111010001","1111111100100010","0000000000100101","0000000011001010","0000000001011110","1111111101010001","1111111100001101","0000000100010001","0000001100010110","0000001001011011","0000000110101000","0000001011100101","0000001000000111","1111111011110101","1111111100110010","0000000101011011","1111111111011111","1111110110011111","1111111011111110","0000000001001001","1111111110000101","0000000000111100","0000000011011010","1111111000111111","1111110101001001","0000000010100010","0000000111101101","1111111110010001","1111111101011111","0000000100100010","0000000011110011","0000000100011010","0000001100001111","0000001011000100","0000000001011111","0000000000000001","0000000001101011","1111111100110011","1111111011001001","1111111110110000","1111111100011111","1111111001110001","0000000000000001","0000000011110100","1111111110111110","1111111110011110","0000000001111001","1111111100001011","1111110101101001","1111111101011111","0000001000110100","0000001000001010","0000000100010011","0000000111101001","0000001001110110","0000000101011110","0000000011001000","0000000100010100","0000000000100010","1111111011000110","1111111111000101","0000000110110010","0000000011100100","1111111001001001","1111110101100000","1111111000001000","1111111001011100","1111111011010111","1111111111100000","0000000000010110","1111111110011000","1111111111001111","0000000000001010","1111111101010111","1111111100111101","0000000000111111","0000000000110010","1111111011000101","1111111001111000","1111111110101010","0000000000101110","1111111110101101","1111111110011111","1111111111000011","1111111011011110","1111110111110100","1111111011110101","0000000011010101","0000000010110111","1111111011100000","1111111001110000","1111111111100001","0000000001111000","1111111110010101","1111111110000001","0000000010001011","0000000010011111","1111111111101101","0000000010010100","0000001000001110","0000000111011011","1111111111110110","1111111010100110","1111111011010010","1111111110000101","1111111111010101","1111111110011010","1111111101000000","1111111101100010","1111111111011110","0000000000001101","0000000001010100","0000000101110001","0000001001000001","0000000101010000","0000000000101010","0000000100111011","0000001100100000","0000001010001101","0000000000101101","1111111110110100","0000000110001011","0000001001000000","0000000001101100","1111111011001101","1111111110010011","0000000100011101","0000000011101111","1111111101010111","1111111010010101","1111111110100010","0000000100010100","0000000100110011","0000000001101111","0000000010010000","0000000101101100","0000000100000111","1111111110000001","1111111100010111","1111111111010100","1111111111001000","1111111100110011","1111111101110101","1111111110100010","1111111011100101","1111111011110001","0000000000111111","0000000010011010","1111111110010101","1111111011101000","1111111010001011","1111110111111001","1111111010010010","0000000000101100","0000000000010111","1111111001011110","1111110111111011","1111111100100010","1111111111000001","0000000000000000","0000000010111111","0000000011000101","1111111101100101","1111111000100101","1111111000100000","1111111011100000","1111111110000111","1111111110000000","1111111101001011","0000000000001101","0000000011101010","1111111111110110","1111111010001011","1111111101111101","0000000110001011","0000000110001000","1111111111100101","1111111100010010","1111111101100110","1111111111000111","1111111101111111","1111111011111001","1111111111001011","0000000111001000","0000000111010011","1111111101111000","1111111001010001","1111111011011111","1111111010101111","1111111110000000","0000001011001010","0000001101001111","1111111100001000","1111110100010110","0000000000000111","0000000110011011","0000000011100000","0000001000011110","0000001010101111","1111111101100011","1111111000000100","0000000110001111","0000001110000000","0000000110011111","0000000011101111","0000000101101100","1111111110111111","1111111000110000","1111111100110111","0000000010011000","0000000101011111","0000001001001100","0000001000100001","0000000101101011","0000001000110100","0000001000001100","1111111100100000","1111110111100000","1111111110110101","1111111110101010","1111110111100110","1111111011110010","0000000010111001","1111111111010001","1111111110110100","0000000110101101","0000000011101111","1111110111000000","1111110101001001","1111111100101101","0000000000001011","0000000001000011","0000000010001111","0000000001110010","0000000011100000","0000000101111101","0000000001110001","1111111101111101","0000000001111100","0000000001111011","1111111011011011","1111111110001011","0000000110010101","0000000011010111","1111111101111100","0000000010000010","0000000100010011","0000000010101011","0000001001100001","0000001110010011","0000000011111100","1111111110100110","0000001001100000","0000001011101101","1111111110100101","1111111011011000","0000000011110100","0000000011101111","1111111110110110","0000000001011001","0000000011001010","0000000000010110","0000000100101000","0000001101011001","0000001011111110","0000000010101000","1111111101111010","1111111111001000","0000000000110011","0000000000101100","1111111111101011","0000000000100100","0000000010100101","0000000000001101","1111111100000101","1111111111111110","0000001000001011","0000000111001101","1111111110110001","1111111010101011","1111111011000111","1111111100001001","0000000001101000","0000000111111100","0000000010001110","1111110100101110","1111110011100010","1111111111101011","0000000110001011","0000000010011111","0000000000110111","0000000010101010","0000000000010110","1111111110000101","0000000001110000","0000000011110001","0000000000010100","0000000000101011","0000000101100100","0000000100001100","1111111101110000","1111111100000101","1111111101100010","1111111101001011","1111111110111100","0000000011010011","0000000100010000","0000000010101101","0000000001100110","1111111101100110","1111111000010001","1111111000101011","1111111100110010","1111111110110100","0000000000100011","0000000010001110","0000000000011100","1111111111011100","0000000010101011","0000000011111000","0000000001101000","0000000001010001","1111111111111010","1111111011100000","1111111100010010","0000000000100101","1111111100110101","1111110110111101","1111111011010110","0000000000011110","1111111011010000","1111110111001111","1111111101010011","0000000011010011","0000000010101011","0000000000000000","1111111101110001","1111111100100110","1111111101011010","1111111110001001","1111111111110010","0000000011110101","0000000010011101","1111111010010100","1111111010111101","0000000101100111","0000000101100110","1111111011011001","1111111101101110","0000001000111010","0000000101111110","1111111010100010","1111111010111110","0000000001000101","1111111101100010","1111110111010110","1111111010001101","0000000001100011","0000000110100100","0000001010010010","0000001011011111","0000000110001001","1111111110000111","1111111011110001","1111111111001001","0000000000101110","1111111110001101","1111111101100001","0000000001000000","0000000010001011","1111111100111111","1111111000100101","1111111101000110","0000000101000010","0000000011111100","1111111010100100","1111110110101111","1111111101000001","0000000011001101","0000000011100100","0000000001101000","1111111101011000","1111110111001001","1111110111011101","1111111110010000","1111111101011010","1111110100110011","1111110110110110","0000000100100111","0000001001000101","1111111111001111","1111111001001001","1111111110000001","0000000001101010","1111111101101000","1111111010000011","1111111100111111","0000000001010011","0000000000110010","1111111110110110","0000000001110110","0000000110000011","0000000011100000","1111111101100010","1111111100111000","1111111111001110","1111111101110111","1111111011111010","1111111101101100","1111111111000111","1111111110110011","0000000001001010","0000000011100000","0000000000010010","1111111100110000","1111111110100110","0000000000000010","1111111111010011","0000000011110100","0000001000111111","0000000010001101","1111110111100110","1111111011001101","0000000110100000","0000000111100110","0000000010101110","0000000100001100","0000000110111100","0000000011110001","0000000001000010","0000000010010000","0000000001101000","1111111110101001","1111111100111010","1111111011000001","1111111001111010","1111111101111101","0000000001111101","1111111110100010","1111111011110110","0000000011001011","0000001010001000","0000000101010110","1111111101101111","1111111101010110","1111111101110101","1111111010101010","1111111011110011","0000000011011100","0000001000001100","0000000101100000","1111111111110100","1111111011011010","1111111010101110","1111111101101101","1111111110101010","1111111010011000","1111110111010111","1111111011001101","0000000000100011","0000000000010011","1111111100001111","1111111011010110","0000000000011001","0000000101111010","0000000100110011","1111111111001001","1111111101000011","1111111111011111","0000000000101101","1111111110101110","1111111011110000","1111111010011101","1111111101110100","0000000011011011","0000000010010110","1111111001100111","1111110100010110","1111110111101001","1111111100000010","1111111100001111","1111111011110100","1111111111010100","0000000110000011","0000001001101000","0000000101101111","0000000000100010","0000000000111001","0000000001101011","1111111110000100","1111111100011101","1111111110111100","1111111110000100","1111111010110101","1111111101010100","0000000010100011","0000000010100001","1111111110001110","1111111001110111","1111110111101110","1111111011000110","0000000001011111","0000000010010001","1111111110010111","1111111110111000","0000000011010110","0000000100100001","0000000010000110","0000000000011000","0000000010100111","0000001001011001","0000001100011100","0000000010101010","1111110111000010","1111111011111111","0000001001100100","0000001000110000","1111111011100000","1111110110101111","1111111101000110","0000000000000001","1111111101000111","1111111110011100","0000000100100010","0000000110110100","0000000100000110","0000000000110101","1111111011101000","1111110100101011","1111110101100001","1111111111110101","0000000100100110","1111111101010101","1111111000110100","1111111111110011","0000000110101000","0000000101000001","0000000001110001","0000000001111111","0000000010011101","0000000000101111","1111111100111011","1111111000000000","1111110101100000","1111110111000110","1111111001010111","1111111010101110","1111111101101010","0000000001101111","0000000011011101","0000000001111010","1111111110010110","1111111011001000","1111111010110110","1111111100100101","1111111101000100","1111111101001010","1111111110101101","1111111111010011","1111111110101101","0000000000000100","0000000000000100","1111111010101000","1111111000000100","1111111111001101","0000000100011011","1111111110001000","1111111000000100","1111111011111001","1111111111100100","1111111100111000","1111111101001101","0000000010001001","0000000001101100","1111111101001011","1111111101110101","1111111111101001","1111111010100100","1111110101100010","1111111001111101","0000000001110100","0000000010010000","1111111100000000","1111111000001011","1111111011001110","1111111111111010","1111111111111111","1111111110111111","0000000010010010","0000000011100011","1111111100100101","1111110110111001","1111111010011010","1111111100111001","1111110111000101","1111110011101011","1111111001101010","0000000000101001","0000000010011111","0000000010000011","0000000001110010","0000000011000101","0000000101101011","0000000011110101","1111111100100001","1111111010010101","0000000010000011","0000001001000011","0000000111101101","0000000011101000","0000000001110110","0000000000000110","1111111101110100","1111111110001111","0000000001000001","0000000000111110","1111111100111001","1111111010110110","1111111101100101","1111111110001011","1111111010100111","1111111100010100","0000000011111111","0000000100101001","1111111101110110","1111111110001000","0000000110000111","0000001000001101","0000000011000111","1111111111110000","1111111111010011","1111111111110101","0000000010011111","0000000011001100","1111111101100011","1111111000011101","1111111010101100","1111111110111101","0000000000100001","0000000011001011","0000000110100100","0000000100000001","1111111100100001","1111111000011101","1111111010011100","1111111110001111","0000000000101111","0000000001000000","1111111111001100","1111111110000101","1111111111011011","1111111111100011","1111111101000100","1111111110011000","0000000100101000","0000000101001001","1111111101011101","1111111011010001","0000000010100011","0000000100100101","1111111101001010","1111111010111010","0000000001010000","0000000010110011","1111111101010100","1111111011110001","1111111110001011","1111111011101101","1111110110110000","1111111000010101","1111111111010011","0000000100000010","0000000100111100","0000000101000001","0000000100100011","0000000010010111","1111111111110111","1111111101111101","1111111010001111","1111110110011001","1111111010001111","0000000100101001","0000001000010011","0000000010100101","0000000000111000","0000000101001110","0000000011000111","1111111100100100","1111111110101010","0000000100001110","0000000001111100","0000000001001001","0000001001111010","0000001101011000","0000000100100011","0000000000010001","0000000101010101","0000000011111100","1111111100010000","1111111110100011","0000001000000011","0000001000010011","0000000000000000","1111111011000111","1111111011011101","1111111101011101","0000000000011010","0000000010000101","0000000000011010","1111111111100100","0000000011101001","0000001001000010","0000001000110010","0000000010000110","1111111100011100","1111111100111001","1111111100110100","1111110111000000","1111110110001011","0000000000110111","0000000111000111","1111111110111110","1111111000011111","1111111100101011","1111111110100100","1111111101011110","0000000110010000","0000001111001100","0000000110110001","1111111010100110","1111111110010011","0000000101100011","0000000000001110","1111111000111011","1111111011100011","0000000001011001","0000000011000110","0000000000111111","1111111100011101","1111111001100100","1111111011100011","1111111110001111","1111111111111010","0000000100110100","0000001000110101","0000000101101000","0000000011010111","0000000111111011","0000000111001011","1111111101010100","1111111011001010","0000000100100001","0000000110010101","1111111011001101","1111110101000000","1111111100000110","0000000011101101","0000000000111000","1111111000110001","1111110110001111","1111111010111111","1111111111001110","1111111111000100","1111111111001111","0000000001111100","0000000011001100","0000000010001000","0000000001000000","1111111111010111","1111111111011111","0000000100100110","0000000110111001","1111111101101001","1111110011100010","1111110111010011","0000000001001000","0000000010000001","1111111101110011","1111111110011010","0000000001010101","0000000001111011","0000000001100110","0000000000001011","1111111110001011","0000000000101101","0000000101010111","0000000011001000","1111111101100010","1111111111011101","0000000100001111","0000000000100110","1111111001010010","1111111000111000","1111111101101011","0000000001110110","0000000011110000","0000000000001100","1111111000011011","1111110111110100","0000000001100011","0000000111101011","0000000010111000","1111111110110010","0000000011011011","0000001000000110","0000000100111000","1111111111001110","1111111110110101","0000000001010001","1111111111001110","1111111010000000","1111111011000011","0000000011001101","0000000110110001","0000000001101011","1111111111001001","0000000100010001","0000000110110010","0000000010110000","0000000001101101","0000000100001010","1111111111011101","1111110111011011","1111111010110101","0000000011110001","1111111111110110","1111110110110000","1111111110010000","0000001100101110","0000000111011111","1111110101101001","1111110011001000","1111111101010100","1111111101100010","1111110110001001","1111111000100000","0000000001001111","0000000010111011","0000000000010111","0000000001101110","0000000011111011","0000000011000001","0000000001110000","1111111111110011","1111111010111101","1111111001101011","0000000001110001","0000001000110110","0000000010011100","1111110111000011","1111110111100011","0000000001001011","0000000100001010","1111111111000110","1111111101000111","0000000000000010","0000000000010011","1111111101001000","1111111100100100","0000000000000111","0000000100001110","0000000110110110","0000000111101101","0000000101011000","0000000000000100","1111111011101101","1111111010111001","1111111100001000","1111111111001010","0000000100001000","0000000101100011","0000000001000010","0000000000110011","0000001000110101","0000001001010110","1111111100101101","1111110111111000","0000000011011010","0000001001111011","0000000011000101","0000000001001011","0000000111101011","0000000111000111","0000000001010010","0000000001100100","0000000001110001","1111111011110110","1111111001111110","1111111110011110","1111111111011111","1111111101110101","1111111110111010","1111111110011010","1111111100110000","0000000000101000","0000000011100100","1111111110001111","1111111011001110","0000000000010101","0000000010001101","0000000000001101","0000000100010000","0000000110110100","1111111110100100","1111111001001110","1111111110110000","1111111111111100","1111111010011000","1111111110010001","0000000111101000","0000000101100111","0000000000000001","0000000100111100","0000001000110111","1111111111100101","1111110110000100","1111111001001001","0000000000111111","0000000011010110","0000000001001100","1111111110110100","1111111101101101","1111111101000110","1111111100100011","1111111110011001","0000000001111100","0000000000000000","1111111001011011","1111111011010101","0000000110111011","0000001011100100","0000000101000100","0000000010000110","0000000101111010","0000000101100101","0000000010000000","0000000010110000","0000000001101111","1111111001111110","1111110111010100","1111111111100100","0000000101001000","0000000000100001","1111111011011001","1111111010111111","1111111001110101","1111110111001100","1111110111100011","1111111011101001","0000000001001110","0000000100010111","0000000001010001","1111111101011001","0000000010110100","0000001100000111","0000001010010011","0000000000010110","1111111101100101","0000000001101111","0000000010100110","0000000001111000","0000000101001010","0000000111010010","0000000100101100","0000000011110100","0000000101110000","0000000010000101","1111111000011101","1111110100010001","1111111010000111","0000000000100111","0000000000001001","1111111101101010","1111111111111110","0000000100010011","0000000101100011","0000000101010001","0000000100111110","0000000001011101","1111111100111101","1111111111001010","0000000101010000","0000000100010111","1111111101101100","1111111100010010","1111111111101101","1111111110011001","1111111010000100","1111111101100110","0000001000010000","0000001100101011","0000000101000011","1111111011000000","1111111001001101","1111111101101011","1111111111101101","1111111101100101","1111111101000110","0000000000010001","0000000001111101","1111111111100000","1111111110000001","0000000000110001","0000000010100100","0000000000010111","0000000000100100","0000000101000001","0000000100000001","1111111100000101","1111111010110001","0000000010111101","0000000110001111","0000000010001000","0000000011110100","0000001010001001","0000001000001001","0000000010101011","0000000110100111","0000001100100001","0000000111101001","1111111111010000","1111111110101001","0000000001101001","0000000001110100","0000000001010000","0000000001011110","0000000000011000","1111111101110100","1111111011001101","1111111011010001","1111111111101010","0000000010100010","1111111110010110","1111111010111011","0000000000001010","0000000101010001","0000000001110001","1111111101101000","1111111111111000","0000000011001100","0000000011111100","0000000010111100","1111111110110111","1111111011110100","0000000000110001","0000000110100001","0000000010101100","1111111100110011","1111111110000101","0000000000000100","1111111111011011","0000000011000100","0000000111011101","0000000100000111","1111111111101110","0000000001110110","0000000011011000","0000000000011000","1111111110110100","1111111110010011","1111111011101101","1111111100101101","0000000011010011","0000000111011011","0000000110000000","0000000010101011","1111111110011101","1111111100010001","0000000000110101","0000000111000101","0000000110101001","0000000010010000","0000000000110000","0000000010000000","0000000011000001","0000000010001101","0000000000001111","0000000001000010","0000000100010110","0000000011110011","0000000001000011","0000000011010101","0000000101011010","0000000000011110","1111111101111011","0000000010010101","0000000010000100","1111111110111001","0000000110101001","0000001110010000","0000000011010001","1111110110001101","1111111011101100","0000000010110111","1111111011000000","1111110101100110","1111111101111011","0000000011100111","0000000000101111","0000000000110110","0000000001010110","1111111001101111","1111110101110100","1111111111110111","0000001000011100","0000000010100100","1111111011010000","1111111110100011","0000000011011100","0000000001011111","1111111110110110","1111111111111000","0000000000010000","1111111110111001","1111111101110101","1111111010110011","1111110110111111","1111111010000000","0000000010100011","0000000101110000","0000000010111011","0000000010011111","0000000011101111","0000000001100001","1111111111011000","1111111111100111","1111111101111011","1111111101011000","0000000011001111","0000000110011110","0000000000011111","1111111101111011","0000000011110110","0000000010101111","1111111000100111","1111110111101011","0000000000001111","0000000001010011","1111111011110011","1111111011011111","1111111101101011","1111111110111111","0000000100001110","0000000110110110","1111111110001100","1111111000000010","0000000000111001","0000001001100000","0000000100110101","1111111110100011","1111111110110000","1111111101110011","1111111010110110","1111111100001101","1111111111100110","0000000000111010","0000000001011001","1111111111100011","1111111010011010","1111111000111101","1111111110010100","0000000010011101","1111111111010100","1111111001001101","1111110111100011","1111111011110100","1111111110101011","1111111011100010","1111111011001110","0000000010101101","0000000101000000","1111111101001010","1111111010110100","0000000000000100","1111111101001001","1111110110100110","1111111100001001","0000000011101101","0000000000101011","1111111111100101","0000000100010001","0000000000000100","1111111001110111","0000000001100000","0000000111111100","1111111111101001","1111111100110101","0000000111001111","0000001000001010","1111111100100111","1111110111111011","1111111010000101","1111111011010010","0000000001011110","0000001000011010","0000000011100100","1111111100110001","0000000000000010","0000000001000100","1111111010111010","1111111100000000","0000000001111100","1111111110101001","1111111001001111","1111111011111000","1111111111010110","0000000010010011","0000001001100011","0000001010110011","0000000010111011","0000000011101010","0000001100000011","0000000111000111","1111111100011101","0000000010000100","0000001010101000","0000000001011010","1111110110100011","1111111011111111","0000000011010011","0000000000001001","1111111100100011","1111111101100001","1111111101011111","1111111110100100","0000000011110111","0000000110101110","0000000011111010","0000000001010000","0000000001000001","0000000000010111","1111111111110000","0000000001000001","0000000010110001","0000000100000001","0000000101100111","0000000110001001","0000000011101001","0000000000010100","1111111110110110","1111111101001110","1111111010111001","1111111101011001","0000000101000101","0000000111101000","0000000001011101","1111111101111111","0000000011010101","0000000111110110","0000000100100111","1111111110100010","1111111011001000","1111111011111010","1111111111011110","1111111111001001","1111111001001001","1111111001100000","0000000101001111","0000001100011000","0000000100101001","1111111010010101","1111110111110011","1111111001000111","1111111011111100","1111111111101111","1111111101110111","1111110111011000","1111110111000000","1111111011100010","1111111010111110","1111111001000101","1111111110100110","0000000101101110","0000000110101011","0000000100010000","0000000000011110","1111111010000100","1111110110100100","1111111010011101","1111111111000100","1111111110100010","1111111100011101","1111111100100111","1111111110110001","0000000001110011","0000000010111001","0000000001001100","0000000010000011","0000000110101000","0000000110010111","1111111111111100","1111111110001111","0000000011110001","0000000101111000","0000000001000100","1111111100110001","1111111100001011","1111111100001000","1111111011100100","1111111100000110","1111111110100100","0000000000100111","1111111101000010","1111110101011001","1111110101010001","1111111110101010","0000000010101000","1111111100110011","1111111100111011","0000000111001100","0000001011000000","0000000011011001","1111111101111011","1111111110111001","1111111110000111","1111111010110010","1111111010111011","1111111110101000","0000000001011000","0000000000101011","1111111110100000","1111111111100000","0000000011001001","0000000010111111","1111111111001110","1111111110001111","1111111110110011","1111111100101100","1111111100100101","0000000000011111","0000000000111110","1111111101110010","1111111110000011","1111111110111100","1111111011011100","1111111010001110","1111111101110010","1111111110000101","1111111100110001","0000000010010011","0000000111100010","0000000010000011","1111111010100011","1111111100000000","0000000000000001","1111111111110000","0000000001001111","0000000111010110","0000001001010101","0000000010110110","1111111100010111","1111111101100010","0000000001101111","0000000001010001","1111111110001010","1111111110011001","0000000000110101","0000000010000110","0000000011001000","0000000010101000","1111111100100111","1111110101000111","1111110100010100","1111110111111010","1111111000011100","1111111000100010","1111111110100010","0000000101101110","0000000100110110","1111111110001110","1111111011110101","1111111110110100","1111111111110010","1111111100111010","1111111010011111","1111111001000011","1111111000110110","1111111110001101","0000000110000101","0000000101111011","0000000000001011","0000000010000010","0000001001010011","0000000111101111","1111111110001100","1111111001100110","1111111100011101","1111111111001000","1111111101100011","1111111010010101","1111111010011011","1111111101110101","1111111101100101","1111111000011100","1111110110110100","1111111001100101","1111111000001001","1111110100010101","1111110111010011","1111111101110111","1111111111100011","1111111110000011","1111111101100000","1111111101011110","1111111110110010","0000000000101001","1111111111010010","1111111110101001","0000000100101111","0000001010000101","0000000110011011","0000000010000001","0000000101010010","0000001000101101","0000000100011110","1111111101001000","1111111001011010","1111111010000000","1111111100010001","1111111110100101","0000000010001100","0000000110000111","0000000011011000","1111111001110110","1111110110101101","1111111110111011","0000000101001111","0000000001111101","1111111100111110","1111111011001001","1111111011011001","0000000000010110","0000000111011101","0000000110101010","1111111111010010","1111111100101010","1111111110111110","1111111111011011","1111111110110101","1111111101001100","1111110111001110","1111110100000000","1111111010110111","0000000000110100","1111111011101000","1111110110110111","1111111100110000","0000000010111000","0000000000111000","1111111111010101","0000000010101001","0000000001110111","1111111010010110","1111110111000011","1111111100110100","0000000000101111","1111111010110110","1111110101000001","1111111010010001","0000000011101000","0000000101101101","0000000010111010","0000000001000111","1111111111000111","1111111110001101","0000000001000000","0000000000110010","1111111010001011","1111110111110010","1111111101001111","0000000000001000","1111111111110010","0000000100010001","0000000111100110","0000000001010100","1111111011000110","1111111110001001","0000000010100010","0000000010010111","0000000010101010","0000000100110110","0000000101111110","0000000110100110","0000000110001001","0000000010101110","1111111111000001","1111111100100101","1111111010010110","1111111101001100","0000000110110001","0000001001010101","1111111101000101","1111110010000011","1111110110010011","0000000000001010","0000000011101001","0000000011011110","0000000011011011","0000000001110001","0000000000101001","0000000010101010","0000000010100110","1111111101101011","1111111011011100","1111111111110111","0000000011010011","0000000010001101","0000000011011001","0000000110101100","0000000010100000","1111111000110100","1111110110100001","1111111011010101","1111111100101000","1111111011101110","1111111110010011","1111111101010000","1111110101110000","1111110110010100","0000000011001111","0000001001010000","1111111111100000","1111110111110010","1111111101111111","0000000110100000","0000000110100111","0000000010001000","1111111011110101","1111110010110100","1111101111110010","1111111010110101","0000000111100100","0000000110000011","1111111110000101","1111111110010000","0000000000111111","1111111110010000","1111111110001010","0000000010101000","0000000000011001","1111111010100110","1111111110000000","0000000011001000","1111111110010110","1111111010011000","1111111111101111","0000000010101110","1111111111100101","0000000000010111","0000000011100001","0000000011010010","0000000101100111","0000001001010010","0000000100100100","1111111111000100","0000000011011100","0000000101010100","1111111101000010","1111111010111001","0000000010100101","0000000010100110","1111111011001111","1111111100010111","0000000010111101","0000000010110010","1111111111000100","1111111110110110","0000000000100001","0000000001011010","0000000000010010","1111111110011100","0000000001110101","0000000111010011","0000000001110001","1111110110000011","1111110111101011","0000000011001001","0000000100111101","1111111111101100","0000000001000111","0000000100101010","0000000010111100","0000000010000110","0000000011110011","0000000001001101","1111111011101100","1111111001000001","1111111010000011","0000000000000011","0000001000010010","0000000111011010","1111111101100001","1111111010011100","0000000000110011","0000000010111001","1111111111000101","1111111110000111","1111111110100110","1111111101011110","1111111111100010","0000000011000101","0000000001000100","1111111110001100","0000000001011001","0000000100111101","0000000100010000","0000000011110001","0000000010101100","1111111100100010","1111110111011110","1111111010010111","1111111110111000","1111111101111001","1111111011100101","1111111101100011","0000000001000111","0000000000001100","1111111010101011","1111111000001100","1111111100011111","0000000000011001","1111111111110010","0000000001100110","0000000110001000","0000000100011110","1111111111110110","0000000001101110","0000000011101101","1111111111001011","1111111111100110","0000001000011101","0000001001001010","1111111110111000","1111111010100101","1111111111000101","1111111111111111","1111111100010101","1111111011110000","0000000000000001","0000000111001010","0000001011101100","0000000111000111","1111111111010100","1111111111011100","0000000010110011","0000000000011101","1111111110000111","1111111111010111","1111111100011000","1111111000101100","0000000000100100","0000001100001101","0000001010101001","0000000001011000","1111111111010101","0000000010010100","0000000010011100","0000000001100111","0000000000111100","1111111101110101","1111111100011100","0000000000011110","0000000011000000","0000000000101100","0000000001010101","0000000101001100","0000000010100010","1111111100010011","1111111101111110","0000000010001101","1111111101010110","1111110111011001","1111111011111111","0000000010011011","0000000000101001","1111111101011111","1111111111001100","0000000000111111","0000000000001101","1111111110000010","1111111010011011","1111111001000110","1111111101000001","1111111111110010","1111111101000011","1111111010100001","1111111010001010","1111111001100010","1111111100011111","0000000010001110","0000000000100110","1111111001011110","1111111001001000","1111111101000000","1111111101000101","1111111111110001","0000000110010000","0000000011101000","1111111010110111","1111111101011101","0000001000001111","0000001011010101","0000001000001011","0000000101010011","1111111111011100","1111111011000011","0000000001100001","0000001001010101","0000000101001100","1111111110001101","1111111111010000","0000000000010000","1111111100110001","1111111110011111","0000000100101111","0000000011001110","1111111011011011","1111111000111110","1111111011101110","1111111101111100","0000000001011111","0000000101110110","0000000011110100","1111111101001110","1111111100010101","0000000000010010","0000000000000010","1111111100101111","1111111100010001","1111111011101111","1111111001010110","1111111100001000","0000000100001000","0000000110111110","0000000010110100","1111111110100010","1111111010010001","1111110110010010","1111111011000101","0000000101101111","0000000101001110","1111111010100001","1111111001000011","0000000000111100","0000000001100000","1111111101000100","0000000000011001","0000000101101011","0000000100000000","0000000010111010","0000000101010110","0000000001100110","1111111001010110","1111111000000011","1111111100000011","1111111101101100","1111111110110110","0000000000111011","1111111111111110","1111111110100100","0000000000111010","0000000010100000","0000000000001110","1111111101110111","1111111011111101","1111111010001000","1111111101110011","0000000101110101","0000000111000100","0000000000001100","1111111100011011","1111111110100111","1111111111000011","1111111100000111","1111111011001110","1111111101100100","1111111111110100","0000000000101110","0000000000111100","0000000000001011","1111111110000000","1111111100110111","1111111111011111","0000000011011111","0000000100000010","0000000010001000","0000000010000001","0000000011001001","0000000010011100","0000000000000110","1111111101110011","1111111101101100","0000000001100101","0000000101100100","0000000011001010","1111111101011000","1111111100010111","1111111110011111","1111111110001001","1111111110001010","0000000000101101","0000000000010001","1111111101110010",
--"0000000001101110","0000000111110100","0000000011000001","1111110111101001","1111110110000010","1111111100111001","1111111101101011","1111111001111110","1111111110110100","0000000111111100","0000000101010101","1111111001110111","1111111000100001","0000000100000000","0000001010101001","0000000100100011","1111111111001000","0000000100101000","0000001011011010","0000000111101001","1111111111001010","1111111110010010","0000000100000010","0000000111110011","0000001000111000","0000001010110110","0000001010111111","0000000101100111","1111111110001010","1111111010011010","1111111100001010","0000000000010010","0000000000011000","1111111011001111","1111111001111010","0000000001100000","0000001000011111","0000000111100010","0000000101000101","0000000100010110","0000000000011101","1111111101110000","0000000011000110","0000000110011100","1111111110100110","1111111000111100","0000000000001001","0000000101111110","1111111111100110","1111111001101000","1111111101110001","0000000011100111","0000000100110011","0000000100011000","0000000010001100","1111111101010011","1111111100001001","0000000010001111","0000000111100101","0000000101100010","0000000001000010","0000000000110111","0000000010101100","0000000001011011","1111111111011011","0000000001000011","0000000001101000","1111111011100111","1111110111101000","1111111111110000","0000001010111111","0000001011010101","0000000110000110","0000000110010101","0000000110001111","1111111101110010","1111110101111111","1111111000111000","1111111111100111","1111111111010101","1111111001111111","1111111000111100","1111111111000011","0000000101010100","0000000100111010","0000000001011100","0000000010100000","0000000101011000","0000000001110110","1111111011000010","1111111011100011","0000000010000101","0000000010100101","1111111100000101","1111111100110001","0000001001001111","0000010000110111","0000001001010011","0000000001101101","0000000101010011","0000000100011001","1111110101111101","1111101110010100","1111111000111100","0000000010011100","1111111111000110","1111111101001111","0000000100011001","0000001001010110","0000000101100101","1111111110100000","1111111011000111","1111111111000001","0000000101000011","0000000100001011","0000000000001000","0000000001100110","0000000010011101","1111111101000000","1111111011110110","0000000001011001","0000000000100111","1111111011101010","1111111111000001","0000000010111101","1111111101011000","1111111010100011","0000000001011110","0000000100100000","0000000000001010","1111111111011001","0000000001110111","0000000001000101","1111111111010100","1111111101000000","1111111000000110","1111110111100111","1111111111000111","0000000100110010","0000000011100011","0000000000011111","1111111101000111","1111111010101100","1111111101101110","0000000001000110","1111111100000110","1111110101011011","1111110111011010","1111111100111000","1111111101011100","1111111011011000","1111111100000011","0000000000010000","0000000100111110","0000000101111101","0000000011111110","0000000011001000","0000000001101000","1111111110101001","0000000000010000","0000000011101010","1111111110110000","1111111000111101","1111111110111011","0000000101100000","0000000001001010","1111111111100010","0000000110010000","0000000100011011","1111111010011100","1111111010110010","0000000001000000","1111111101011111","1111111000110001","1111111111000001","0000000110010101","0000000100110101","1111111111100110","1111111011010010","1111111001000100","1111111011001111","1111111101101111","1111111010011100","1111110111011101","1111111101100011","0000000110111111","0000001000100001","0000000010100111","1111111110110001","0000000000110011","0000000010000011","1111111101111100","1111111011111001","0000000001000110","0000000011110000","1111111110000111","1111111100011001","0000000101001111","0000001100000110","0000001001011001","0000000101101100","0000000110000011","0000000101110000","0000000011110101","0000000011101011","0000000011100001","1111111111001111","1111111001101001","1111111011000000","0000000011100110","0000000111011111","0000000001101000","1111111110111000","0000000100111101","0000000101111101","1111111111100001","0000000010110010","0000001101011001","0000001001100100","1111111100001000","1111111100011010","0000000101011011","0000000100001011","1111111110111010","0000000001000111","0000000010010110","1111111110111000","0000000000110000","0000000101111011","0000000100010001","0000000000000001","1111111111111000","0000000000100000","0000000010010110","0000000110101111","0000000100100111","1111111011111001","1111111011111100","0000000011101011","0000000010010101","1111111100000000","1111111110100000","0000000000100001","1111111001101011","1111111011001110","0000001001111010","0000001110010010","0000000011101000","1111111111110010","0000000100101101","0000000010000100","1111111011111010","1111111110011100","0000000001100111","1111111101110100","1111111101100001","0000000100000001","0000000101101010","0000000000111001","1111111110101111","1111111111010101","1111111110100101","1111111110010110","1111111110100001","1111111011100111","1111110111110001","1111110110100101","1111111000001111","1111111110010111","0000000110110010","0000000110101011","1111111101011101","1111111010010000","1111111111110000","1111111111110010","1111111010100101","1111111101011001","0000000100010010","0000000100000111","0000000011001101","0000000111000011","0000000101101011","1111111110111011","1111111111101101","0000000110000101","0000000111110001","0000000111110111","0000000111011010","1111111110010101","1111110101011100","1111111100101001","0000000111100001","0000000010111001","1111111010101010","1111111110010110","0000000010110100","1111111111010000","1111111110010111","0000000011000110","0000000100100011","0000000010110000","0000000000110101","1111111011100001","1111110101111110","1111111000010010","1111111110001110","1111111110010010","1111111001101000","1111110111110101","1111111101100100","0000000111101111","0000001010100111","0000000001111010","1111111010111001","1111111100111010","1111111101110101","1111111100101010","0000000010101111","0000000110111110","1111111101010001","1111110101111011","1111111111000001","0000000101101111","1111111101101100","1111111001101000","0000000001101100","0000000011101110","1111111011000011","1111111000011110","0000000000100010","0000000110101110","0000000101000010","0000000000111011","1111111111010001","1111111111010111","1111111111111000","0000000001111110","0000000011111000","1111111111111010","1111111001000101","1111111011001110","0000000101100100","0000001001110111","0000000101011010","0000000010000001","0000000001010001","1111111110111100","1111111100110001","1111111100011011","1111111100011000","1111111101101011","1111111111000110","1111111100110100","1111111011011110","0000000000010111","0000000100000110","0000000000101110","1111111100110010","1111111011001110","1111111001011011","1111111100010101","0000000101000010","0000000111111100","0000000010100001","1111111111101011","0000000001001110","0000000010101000","0000000111001110","0000001101100111","0000001011011010","0000000010010100","1111111110010100","0000000000100100","0000000011100110","0000000101111111","0000000101100001","0000000010001110","0000000010100011","0000000100110000","0000000000000000","1111111001100101","1111111100100000","0000000011001011","0000000101011100","0000001000000111","0000001010110100","0000000100100011","1111111010101010","1111111010101101","0000000001101010","0000000100110110","0000000101001101","0000000110000101","0000000011100011","1111111101001110","1111111010001111","1111111101111101","0000000010101011","0000000001000110","1111111001010100","1111110100011101","1111111001111100","0000000100100010","0000001000111011","0000000100110011","1111111111011111","1111111101011001","1111111100111000","1111111110100000","0000000011101010","0000000101100001","1111111111001001","1111111011010101","0000000001100101","0000000011110000","1111111010010010","1111110111011101","0000000010001101","0000000110100011","1111111111101101","1111111111010101","0000000100110100","0000000010001000","1111111101101010","0000000000111110","0000000011001001","0000000001010110","0000000011010010","0000000010100000","1111111001000001","1111110110000101","1111111111110100","0000000100101001","1111111111000101","1111111011111011","1111111101011101","1111111111001011","0000000010111101","0000000100000010","1111111100110010","1111111001101010","0000000010100000","0000000110000011","1111111011000001","1111110011001100","1111111001000000","0000000000101101","0000000010111010","0000000100000010","0000000100101011","0000000010000001","1111111110000111","1111111101100010","0000000010010111","0000001000010111","0000000111000100","1111111111010011","1111111101010000","0000000011011110","0000000101100100","1111111111010011","1111111011011001","1111111110100110","0000000001000010","1111111101111011","1111111001011100","1111111000010100","1111111011100111","0000000001010101","0000000100001100","0000000001010010","1111111110011111","0000000010001110","0000000110101011","0000000010011110","1111111010101110","1111111011010010","0000000001101010","0000000010100101","1111111110011000","1111111101000101","1111111111010011","0000000001000101","0000000001100111","0000000000001110","1111111100111110","1111111100000011","1111111111000111","0000000001110011","0000000001100110","0000000000001011","1111111111000110","0000000000000110","0000000010101001","0000000000111010","1111111010111110","1111111011001011","0000000010000100","0000000001100100","1111111000001111","1111110101101011","1111111100110001","0000000000100011","1111111111001111","0000000010001010","0000000111111101","0000001000011101","0000000100011011","0000000000001010","1111111100000011","1111111001100101","1111111010100100","1111111011101000","1111111010000110","1111111001000011","1111111010110000","1111111101111001","0000000000111110","0000000000111011","1111111011011011","1111110111001111","1111111011111010","0000000001001110","1111111100011011","1111110110101101","1111111100111011","0000000101001110","0000000000110101","1111110111110011","1111111001000100","0000000001101000","0000000110010101","0000000100101011","0000000000010000","1111111110100111","0000000011111010","0000001010100100","0000001001110010","0000000100111000","0000000011001000","0000000001101001","1111111110100100","1111111111001111","1111111111101010","1111111000000111","1111110011111010","1111111111010001","0000001011010100","0000000111110101","1111111111111110","0000000000010100","0000000010000100","0000000001101010","0000000011011010","0000000000000111","1111110100001011","1111110010010100","0000000010111101","0000001110101000","0000000110110000","1111111101000111","1111111110001111","1111111110111000","1111111010100101","1111111011111001","0000000010001110","0000000010101011","1111111111000110","0000000000100000","0000000100001010","0000000010011100","1111111101111100","1111111101011111","0000000000101010","0000000010100010","0000000000110001","1111111101001101","1111111011111011","1111111110100010","0000000001010011","0000000000011010","1111111101001000","1111111010011011","1111111001001000","1111111001100010","1111111011100010","1111111101010101","1111111101010110","1111111100011001","1111111101000111","0000000001011100","0000000110001100","0000000101000110","0000000000010111","0000000001011000","0000000110000001","0000000010111110","1111111100000011","1111111110000100","0000000011110101","0000000001111100","0000000000011000","0000000111001101","0000001010100010","0000000100101110","0000000010111111","0000000110110110","0000000011000011","1111111010011110","1111111001111110","1111111101001010","1111111011010011","1111111010011111","1111111101111110","1111111100111100","1111110111101100","1111111000111110","0000000000001011","0000000011011000","0000000001111100","0000000001000101","1111111111111000","1111111100110101","1111111011111100","1111111101101000","1111111100101010","1111111010001100","1111111101010100","0000000011111100","0000000110000100","0000000101100000","0000000110110100","0000000100100111","1111111101110110","1111111101011101","0000000010110101","0000000000110101","1111111011000101","1111111110010011","0000000001101101","1111111010011011","1111110110100011","1111111111001000","0000000100000011","1111111111011100","1111111110101101","0000000000011111","1111111010100111","1111110111010101","1111111111111101","0000000101001110","1111111101011010","1111110111010001","1111111100010101","0000000011011101","0000000101110010","0000000101001000","0000000010110001","1111111111110101","1111111110111011","1111111111101100","0000000000001100","0000000000110100","0000000010111000","0000000101110100","0000000110001111","0000000001100111","1111111011111100","1111111010111111","1111111100110001","1111111101110110","0000000000110001","0000000100110010","0000000100011111","0000000010101101","0000000100010111","0000000011110010","1111111111011010","0000000000101001","0000000101000010","0000000000111110","1111111100011001","0000000011100101","0000000111100111","1111111010110010","1111110001001110","1111111011000111","0000000110010001","0000000100111111","0000000100100010","0000001001100000","0000000110101100","1111111101100011","1111111100100010","0000000010000011","0000000010110100","1111111111001111","1111111100100001","1111111010100101","1111111010100101","1111111110011010","0000000001111100","0000000001101000","1111111111111010","1111111110000011","1111111100000100","1111111110011100","0000000110101010","0000001011101100","0000000101111110","1111111100000010","1111111010000000","0000000000001001","0000000010000011","1111111001110101","1111110011100111","1111111001111101","0000000010000111","0000000000000011","1111111101001010","0000000011010101","0000001001011011","0000001000101100","0000000111010110","0000000101010101","1111111111111110","0000000000011101","0000000111011010","0000000101001100","1111111100001001","1111111110101101","0000000110010001","0000000001001100","1111111010111000","0000000001111010","0000000111110111","0000000010111111","0000000000010100","0000000001110001","1111111110010011","1111111101010010","0000000100000010","0000000100100001","1111111100100001","1111111011000000","1111111110001010","1111111011101101","1111111011100111","0000000011010111","0000000110101001","0000000010111010","0000000001110101","0000000001101101","1111111111011100","0000000001110010","0000000011100111","1111111010011100","1111110011111000","1111111101111001","0000000110101111","0000000000100101","1111111100111101","0000000100010010","0000000101101100","1111111110111110","1111111110011011","1111111111101111","1111111000111001","1111110101000001","1111111100010100","0000000001001100","1111111101001110","1111111011110000","1111111111000000","1111111101110110","1111111010011100","1111111100101111","0000000000000000","1111111100000010","1111110101001000","1111110100110000","1111111010110101","1111111111010100","1111111110101001","1111111101111000","0000000001000000","0000000100001001","0000000011010000","0000000000000010","1111111100001100","1111111001000100","1111111011000110","0000000001010001","0000000011001010","1111111111111100","1111111110011101","1111111101101011","1111111011101010","1111111111110011","0000000111100111","0000000100000010","1111111001111100","1111111101010100","0000000111101011","0000000100001000","1111111011000001","1111111111101110","0000001001001001","0000000110011010","1111111101101001","1111111010111010","1111111101100101","0000000000000001","1111111101000101","1111110110100011","1111111000111110","0000000101000001","0000000110011110","1111111001011010","1111110100000100","1111111010101100","1111111011100010","1111111000101110","1111111111010010","0000000101010000","0000000000100001","1111111101100111","0000000001000101","1111111111111100","1111111110011110","0000000100111011","0000000110010110","1111111100101000","1111111000110000","1111111101011100","1111111010110100","1111110101000111","1111111011110101","0000000110100000","0000000101100011","1111111110010110","1111111010111110","1111111001101101","1111111000010010","1111111001101010","1111111111110111","0000001000001110","0000001010011000","0000000011001111","1111111110110011","0000000011111000","0000000110010001","0000000010011110","0000000101100100","0000001011011010","0000000101000110","1111111110011001","0000000110101110","0000001100101111","0000000010001110","1111111001001111","1111111100010100","1111111101110111","1111111011001011","1111111101011101","0000000000110111","1111111111010100","1111111100110011","1111111010110011","1111111001101101","1111111110000000","0000000001111101","1111111100001001","1111110101110001","1111111010001100","0000000000001011","1111111110110000","1111111100110100","1111111101110100","1111111110000001","1111111110111010","0000000001001001","0000000001100101","0000000010110111","0000000101100111","0000000010110100","1111111101011011","1111111110111111","0000000001010011","1111111100010010","1111111001111101","1111111111101011","0000000001101001","1111111110000000","1111111110110001","0000000000000100","1111111010101100","1111111000011011","0000000000001101","0000000110111100","0000000100110101","1111111111011101","1111111101000100","0000000001011100","0000001011010001","0000001101110010","0000000010000101","1111111000010001","1111111101101010","0000000101010111","0000000011010001","0000000000101100","0000000010101001","0000000000010001","1111111101100010","0000000101110101","0000001100110101","0000000001101001","1111110011111111","1111111000111111","0000000100001010","0000000100000000","0000000010000001","0000000101110110","0000000011111100","1111111100010000","1111111101000010","0000000011011010","0000000011011011","0000000010001010","0000000101001100","0000000010010100","1111110111110011","1111110100100000","1111111011111000","0000000000011101","1111111100010111","1111110111111100","1111111001110011","1111111110010101","1111111111110000","0000000000100111","0000000101111010","0000001000100111","0000000000110010","1111111010010111","0000000001101001","0000001001100111","0000000110000100","0000000011001000","0000000110110001","0000000011011111","1111111010011000","1111111010011000","1111111110100111","1111111011011000","1111111001011001","1111111110100011","1111111110110001","1111111010001111","1111111110000111","0000000011111011","1111111110101101","1111111001111111","0000000001110101","0000001000000100","0000000001010110","1111111010101101","1111111110000101","0000000010110110","0000000001111010","1111111110100101","1111111101001010","0000000000011101","0000000111000100","0000000111101001","1111111110001010","1111110110101001","1111111010111110","0000000010110000","0000000011001100","1111111110101100","1111111011110001","1111111011111000","1111111110010110","0000000000110110","0000000000001111","1111111110010101","1111111111001111","0000000010011101","0000000101101001","0000000111001101","0000000100010011","1111111110101100","1111111101101110","0000000000101110","0000000001101000","0000000100010101","0000001011100000","0000001001110110","1111111011000100","1111110011010111","1111111011111110","0000000010101100","1111111101110001","1111111001100100","1111111100110111","0000000001010110","0000000001110101","1111111101000110","1111110111111001","1111111011110001","0000000100101111","0000000011000011","1111111001000011","1111111000000111","1111111110111010","1111111111000010","1111111001111101","1111111001111011","1111111101110001","1111111111011110","1111111110001100","1111111100110010","1111111111001000","0000000011100011","0000000010001111","1111111100010000","1111111011111101","0000000000100100","0000000000100011","1111111101001100","1111111100011111","1111111011111010","1111111001110001","1111111010001111","1111111110000110","0000000011111011","0000001001011000","0000000110101110","1111111100010111","1111111001111100","0000000010101001","0000000110010110","0000000011111100","0000000111111011","0000001010001000","1111111110100001","1111110101100100","1111111100110010","0000000010111010","1111111110101001","1111111111100001","0000000100100100","1111111011011101","1111101101001001","1111110001100011","0000000000101100","0000000011001110","1111111101010000","1111111101100010","1111111110010000","1111111000111100","1111111001111000","0000000101001101","0000001001110001","0000000001110011","1111111110100011","0000000101111011","0000000111110011","1111111111011000","1111111100101111","0000000101110101","0000001011110110","0000000101101011","1111111101000001","1111111100010110","0000000000010110","0000000000110110","1111111101101011","1111111011101111","1111111011010001","1111111010010110","1111111100011110","0000000011011100","0000000110111100","0000000000101110","1111111001001111","1111111010110001","0000000001101110","0000000100010011","0000000000100000","1111111100010110","1111111101011111","0000000010010100","0000000011111010","0000000000111100","0000000000000111","0000000100000110","0000000111010000","0000000101001111","1111111111100101","1111111010011100","1111111010001101","1111111110110100","0000000010100001","0000000011010001","0000000011101110","0000000001001110","1111111011000000","1111111011000111","0000000010011110","0000000001001110","1111110111011111","1111111001001101","0000000100000011","0000000010101111","1111111011010100","0000000001000100","0000000111110001","1111111110010000","1111110101111000","1111111110010010","0000000101101110","0000000000001010","1111111011110100","1111111110010100","1111111111011101","0000000010010110","0000001001110100","0000001000110100","1111111100010111","1111110101100100","1111111010010110","1111111110110000","1111111111000011","0000000001001000","0000000011100001","0000000010000111","1111111111110010","0000000000000001","0000000001000100","1111111111000100","1111111001100001","1111110111100111","1111111111001100","0000000110011101","0000000001111011","1111111100000001","0000000001110011","0000000111000011","1111111111001011","1111111000100111","1111111110000001","1111111111101000","1111110110111110","1111110111001111","0000000101100010","0000001100111100","0000000100100111","1111111010100111","1111111000001010","1111111001111001","1111111101000011","0000000000100001","0000000010011010","0000000011011001","0000000011000001","1111111111011110","1111111110001010","0000000011111010","0000000111010001","0000000001011110","1111111110001010","0000000001111101","1111111110110000","1111110101001100","1111110111011011","0000000000011111","1111111101000011","1111110110100111","1111111110100101","0000000110100000","0000000000110110","1111111110011001","0000000101001111","0000000011000111","1111111010001100","1111111100100100","0000000001110001","1111111011101000","1111111000010000","0000000001101010","0000000111100100","0000000010011001","1111111100001110","1111110111010010","1111110100000100","1111111010000010","0000000001101111","1111111100011010","1111110100011101","1111111010010101","0000000010110100","0000000000000000","1111111100000101","1111111111110011","0000000010101110","0000000001010110","0000000001000111","0000000000111010","1111111101111100","1111111100110100","0000000000100010","0000000100011101","0000000011001011","1111111110000000","1111111101110010","0000000110100011","0000001100111001","0000000110011010","1111111100111011","1111111101000100","0000000001011011","0000000001011111","1111111111001110","1111111011101101","1111110110011000","1111110101110001","1111111011100110","1111111111001111","1111111111101111","0000000011001111","0000000101000101","0000000000011101","1111111110100011","0000000010111111","0000000011101110","0000000001000111","0000000100010111","0000000111000001","1111111111101001","1111111001011011","1111111110110000","0000000100111111","0000000011000111","1111111111111010","1111111111110000","1111111110011011","1111111011011010","1111111010000010","1111111011110101","0000000000111000","0000000101011000","0000000100001110","0000000000011000","1111111111101001","0000000000011011","0000000001010000","0000000011110101","0000000011000101","1111111100100010","1111111100101001","0000000111011101","0000001011100001","0000000011101000","0000000000111000","0000000101110100","0000000100100000","0000000000001111","0000000010101101","0000000001110011","1111111000000110","1111110110101101","0000000010001010","0000000111010100","0000000000000011","1111111001011001","1111110111110110","1111111000111111","1111111111111100","0000001000011010","0000000110101101","1111111101101101","1111111001111111","1111111011100010","1111111011010010","1111111010001000","1111111011010011","1111111110000000","0000000000011111","0000000000000110","1111111101010111","1111111111101101","0000000110111001","0000000110000011","1111111101000001","1111111011110100","0000000001110011","1111111110101110","1111110110001100","1111111000011000","0000000000011101","0000000001100100","1111111111101110","1111111111100000","1111111011010111","1111110111011000","1111111100010001","0000000000110011","1111111010110001","1111110101111110","1111111100111001","0000000011111101","0000000001001100","1111111101010101","0000000001001101","0000000111100000","0000000110011001","1111111101101101","1111111000100101","1111111110010100","0000000100110011","0000000000100110","1111111001110101","1111111011001111","1111111100111101","1111110111111010","1111110110110011","1111111110101111","0000000011010001","1111111110111101","1111111011001010","1111111011100010","1111111100001110","1111111111001111","0000000110011111","0000001011010110","0000001001000010","0000000011101010","0000000000001111","0000000000100101","0000000100110100","0000001001011110","0000001000111001","0000000011000100","1111111111000000","0000000010000000","0000000111100101","0000000110001101","1111111101010100","1111110111111011","1111111011110010","0000000001000111","0000000000110110","1111111101101011","1111111011111010","1111111110000010","0000000100001110","0000000101111001","1111111011111001","1111110011100111","1111111100110111","0000001010011011","0000000110110011","1111111011001000","1111111011101000","0000000001110011","1111111110011110","1111111001010011","1111111101111111","0000000011010110","1111111111010101","1111111011101010","0000000001000100","0000000100000111","1111111011001001","1111110011000100","1111111001000110","0000000010100110","0000000001100101","1111111100110111","1111111101101101","1111111101011011","1111111000111110","1111111010010111","0000000001000011","0000000000101011","1111111100000010","1111111111011111","0000000101011101","0000000010011011","1111111110000100","0000000010111001","0000001000110100","0000000110110011","0000000010110000","0000000001110111","0000000001011010","0000000010100010","0000000110000110","0000000011111101","1111111011000100","1111111001100101","0000000011010010","0000001000000101","0000000001100010","1111111100111000","1111111111001100","1111111110110011","1111111011001110","1111111101101011","0000000011110100","0000000100001100","0000000001000110","0000000011000000","0000001000011100","0000001001100001","0000000011100101","1111111011100110","1111111001000101","1111111101111110","0000000010111101","0000000001010000","1111111101000000","1111111101000011","1111111111101010","0000000001011001","0000000100011110","0000000111100000","0000000010111100","1111111000111001","1111110110001001","1111111100011100","1111111111110011","1111111101011010","1111111101100100","1111111111011000","1111111100010010","1111111001010010","1111111101010110","0000000010010000","0000000000100010","1111111011011010","1111110111101110","1111110111110101","1111111101101000","0000000100011100","0000000101010011","0000000011111100","0000000100001111","1111111110100110","1111110100100100","1111110101100110","1111111111010010","0000000000000010","1111111100010000","0000000001100101","0000000011101010","1111111000000011","1111110100000001","0000000010010101","0000001010010110","0000000000110010","1111111001110101","1111111100100000","1111111100110110","1111111101101110","0000000101000110","0000000100100000","1111110110101001","1111110000101001","1111111010010001","1111111111111011","1111111010011010","1111111000000001","1111111011011110","1111111011000000","1111111001001111","1111111101011100","0000000000110010","1111111100101111","1111111010100000","0000000000111010","0000000110001101","0000000001110110","1111111011100011","1111111100100001","0000000000010100","1111111111101110","1111111110000111","0000000000000101","0000000000011100","1111111100001000","1111111010111111","0000000001001100","0000000111011000","0000001000000110","0000000100010100","1111111100100110","1111110110101010","1111111100000001","0000000101101010","0000000010010100","1111111000001001","1111111100010100","0000001010000000","0000001011101011","0000000011011110","0000000001111001","0000000101010111","0000000011110110","0000000000001110","1111111111011011","1111111101110110","1111111010100110","1111111010111000","1111111111011101","0000000011010101","0000000011111000","0000000011000000","0000000010101010","0000000010110110","0000000011100000","0000000011110011","1111111111111001","1111110111101101","1111110101010100","1111111110000010","0000000101101100","0000000011010101","0000000000010000","0000000000110111","1111111100001010","1111110110011111","1111111100101111","0000000101001110","0000000001101111","1111111111011110","0000001001000001","0000001010111110","1111111101000100","1111110110001110","1111111101111000","0000000000101010","1111111100011000","1111111111000111","0000000011100111","0000000000010101","1111111111001011","0000000011100111","0000000000111111","1111111010111101","0000000000100101","0000001001000111","0000000101000101","1111111110011011","0000000000111000","0000000011011110","0000000010001001","0000000100100100","0000000110000001","1111111111101110","1111111100011001","0000000000100101","0000000000000111","1111111100011001","0000000001101101","0000000110100101","1111111110000011","1111110110100101","1111111101010100","0000000100101111","0000000011100010","0000000010110010","0000000011000111","1111111110000010","1111111010110111","0000000000001001","0000000100000110","0000000000001001","1111111010111100","1111111001000110","1111111001011000","1111111010100010","1111111010100100","1111111011101010","0000000011010101","0000001010011001","0000000101001111","1111111110001110","0000000101000101","0000001101001011","0000000100101111","1111111000101000","1111111011000110","0000000011110101","0000000101010000","0000000001111011","1111111111001010","1111111100111111","1111111100010001","1111111101001000","1111111110111010","0000000011000001","0000000110000110","0000000011001100","0000000000110010","0000000100101100","0000000100011110","1111111011001110","1111110111111110","0000000000010011","0000000110001110","0000000100100001","0000000001011110","1111111100101101","1111111000111110","1111111111100111","0000001001010000","0000000110001101","1111111101010001","1111111100000010","1111111011101111","1111110111010000","1111111010000011","0000000011011101","0000000010101010","1111110111110111","1111110100000000","1111111010101100","0000000001010110","0000000010001111","1111111111011001","1111111100101110","1111111101011010","0000000000110001","0000000010011110","1111111111100101","1111111010011011","1111111000110100","1111111100010111","1111111111000001","1111111101101101","1111111110001101","0000000001111111","0000000010101111","0000000000000100","1111111101101010","1111111001111111","1111111000101001","0000000000111011","0000001000101011","0000000010010010","1111111010110010","0000000001100110","0000001000001100","0000000000110001","1111111000101100","1111111001011110","1111111010111101","1111111100011010","0000000000111110","0000000000100111","1111111011110000","1111111111000011","0000000110101000","0000000101010001","0000000000111111","0000000010011100","0000000001110010","1111111110000100","0000000010001010","0000001001010001","0000000111010111","0000000011000111","0000000100011100","0000000011010100","1111111111000010","0000000010110001","0000001010010010","0000000111111111","0000000000100001","0000000000000100","0000000011100010","0000000011000110","1111111111110110","1111111100100111","1111111010010100","1111111010111100","1111111101101011","0000000000100001","0000000101100000","0000001010100111","0000000111010110","1111111101101000","1111111010111010","0000000000100001","0000000011000101","0000000001101110","0000000100011011","0000001000100011","0000000110011011","0000000000111100","1111111111000010","0000000000011010","0000000010000111","0000000010111000","0000000001011011","1111111111010111","0000000001001011","0000000101011000","0000000100100111","1111111110110110","1111111100101101","0000000000001100","0000000000001010","1111111001001101","1111110110101000","1111111111100110","0000000111110011","0000000010110111","1111111010011111","1111111101001001","0000000101001010","0000000101100100","1111111111111010","1111111100010001","1111111100001000","1111111110100110","0000000010100000","0000000011111010","0000000001111011","1111111111101000","1111111101010011","1111111100010110","0000000000110111","0000000100111100","1111111111000010","1111110111010111","1111111010101100","0000000000101011","1111111110000001","1111111010100110","1111111101000101","1111111110100101","1111111110001010","0000000000010011","1111111111111001","1111111011101010","1111111101100111","0000000100101010","0000000100110010","1111111111110101","1111111111001010","0000000000111000","0000000001110111","0000000100110001","0000000110010110","0000000001110010","1111111100010101","1111111010111111","1111111011111011","1111111110111000","0000000010010111","0000000000000110","1111111001001101","1111110110010110","1111111001001100","1111111110110001","0000000110000000","0000001001010000","0000000101001011","0000000010111110","0000000110000100","0000000011100000","1111111100101011","1111111111111010","0000001000000010","0000000101101001","0000000000001100","0000000100000110","0000000111000110","0000000001000100","1111111110001100","0000000010100100","0000000001110011","1111111011001100","1111111001110001","1111111100110111","1111111101001011","1111111011111110","1111111100011001","1111111101111010","0000000001101110","0000000110001000","0000000011100010","1111111010011111","1111110101110010","1111111000100110","1111111011100101","1111111011000000","1111111001010111","1111111010000000","1111111111011110","0000000101111000","0000000100000110","1111111101011000","1111111111000010","0000000101100001","0000000010011111","1111111101000110","0000000011100000","0000001001000101","1111111111010001","1111110111000011","1111111111011110","0000000111100110","0000000011000111","0000000000010111","0000000101010000","0000000100110001","1111111101101110","1111111011111101","0000000000111011","0000000110101001","0000001001011001","0000000011101010","1111110110101001","1111110001000001","1111110111101000","1111111100011000","1111111010100001","1111111101000100","0000000010100010","1111111110110100","1111110110110001","1111111000011001","0000000001100100","0000000111001010","0000000110010000","0000000000101110","1111111010101011","1111111100000101","0000000101010110","0000001010110110","0000000110101001","1111111111110111","1111111100110010","1111111101001100","1111111110100011","1111111100110000","1111111000100001","1111111010010100","0000000010000000","0000000010110011","1111111011111000","1111111010111000","1111111111100111","1111111110110110","1111111100001001","1111111110101010","1111111110001100","1111110111100110","1111110111000100","1111111101111001","0000000000101001","1111111111101000","0000000000011001","1111111110110101","1111111011100001","1111111101011000","1111111110110011","1111111010000001","1111111010111101","0000000100010100","0000000011100100","1111111000000000","1111110111111010","0000000011011111","0000000110001100","0000000001101011","0000000100111100","0000001000110101","0000000001100100","1111111010010110","1111111110010000","0000000011000100","0000000000010011","1111111100110001","1111111011101011","1111111000111110","1111110111111000","1111111100010111","1111111111011111","1111111101001101","1111111100100111","1111111111001111","1111111110100110","1111111101110001","0000000010100101","0000000101000011","1111111111101000","1111111100110101","0000000000011100","0000000000010110","1111111101110011","0000000010100010","0000001000100111","0000000110111100","0000000100000110","0000000100000100","0000000000100101","1111111101000011","0000000000000101","0000000010000110","1111111110111110","1111111111001001","0000000000011111","1111111010100001","1111110101110101","1111111010111110","1111111111001000","1111111100100010","1111111100101000","0000000000011101","0000000010110110","0000000110110110","0000001001111011","0000000011101011","1111111100100000","0000000000111010","0000001000000000","0000000111010010","0000000100010001","0000000001101101","1111111110000011","0000000000100101","0000001000110110","0000001000011011","1111111111100101","1111111100001001","1111111101010110","1111111100110010","1111111110101101","0000000001000101","1111111101101101","1111111110100011","0000001000000011","0000000111111100","1111111011011010","1111111000101010","0000000001000001","0000000010011000","0000000001000011","0000000111000001","0000000110100101","1111111011011000","1111111001000110","1111111111111010","1111111100111110","1111110111010101","1111111111110111","0000001001010000","0000000100101001","0000000000111100","0000000111000100","0000000111010110","1111111111111000","0000000001010011","0000001000011101","0000000101001010","1111111110000010","0000000001011111","0000000110010001","1111111111001001","1111110110101000","1111111011100000","0000000111000111","0000001010000000","0000000010110000","1111111100000000","1111111011100000","1111111100000100","1111111001110011","1111111010100011","0000000001001001","0000000100010011","0000000000001001","1111111111010000","0000000100101101","0000000101010001","1111111111110000","1111111110111101","0000000001110000","1111111111110011","1111111110000010","0000000011000011","0000000111100000","0000000101001110","0000000000111101","1111111100111101","1111110111110000","1111110101011001","1111111001010101","1111111111101001","0000000011011010","0000000001110101","1111111100000000","1111111001111000","1111111110011111","0000000000010010","1111111100110000","1111111110111110","0000000101001000","0000000010000010","1111111100110100","0000000100001110","0000001011111100","0000000011100000","1111111000101001","1111111011110101","0000000011101000","0000000101011101","0000000101100011","0000000011110101","1111111101011001","1111111010110000","0000000000001011","0000000010110001","1111111111000010","1111111111010100","0000000100110000","0000000101010101","0000000000001100","1111111100101100","1111111100110011","1111111111000010","0000000011000000","0000000100010110","1111111101011110","1111110011100011","1111110011101101","1111111110111110","0000000101010000","1111111101000111","1111110100010110","1111111001001010","0000000010010010","0000000010001010","1111111111000111","0000000010011111","0000000101111000","0000000011110011","0000000010100001","0000000010111000","1111111111001010","1111111011110100","1111111111001100","0000000001101011","1111111101001010","1111111011001001","0000000001011010","0000000110011100","0000000100011110","0000000010001101","0000000010100001","0000000000000011","1111111011001000","1111111010101111","1111111111111100","0000000101001111","0000000111011001","0000000101000100","1111111011111000","1111110001001000","1111110011000000","0000000010001110","0000001001101001","1111111110011000","1111110011111010","1111111010110111","0000000101111010","0000000101101011","0000000001101100","0000000010100101","0000000001011011","1111111010110111","1111110111011110","1111111010110101","0000000000000010","0000000101100110","0000001011110111","0000001110110011","0000001100010001","0000000111011001","0000000001110100","1111111011100000","1111111000010001","1111111011101011","0000000001110101","0000000011101000","1111111111010101","1111111001110101","1111111001010101","1111111110011101","0000000010011011","0000000000101111","1111111111001000","0000000010101111","0000000011100110","1111111010001110","1111110010010011","1111111010100110","0000001000111101","0000000111110011","1111111010110000","1111111000110111","0000000100101100","0000001010011000","0000000100011001","0000000000010100","0000000000100011","1111111100010111","1111111000111001","1111111110100001","0000000010011001","1111111011111000","1111111000010001","1111111110000001","1111111111011111","1111111011101011","1111111111100011","0000000100010101","1111111100101010","1111110101001000","1111111011101010","0000000011010101","0000000001001011","1111111110000010","1111111101001100","1111111001111110","1111111001111000","0000000000001001","0000000011110101","0000000011111101","0000000110101110","0000000110111000","0000000000100001","1111111101110000","0000000000110111","1111111111110101","1111111100001100","1111111110110010","0000000011111000","0000000101000111","0000000101000001","0000000101000000","0000000011111011","0000000011110100","0000000011100101","0000000001001011","0000000001011010","0000000100101001","0000000010100100","1111111101010101","1111111110011100","0000000000011011","1111111011110011","1111111010100100","0000000010000001","0000000101001000","1111111111010111","1111111011111000","1111111101101010","1111111110111110","1111111111111011","0000000000101011","1111111101110101","1111111010011111","1111111100011011","0000000001001111","0000000010100101","1111111100111110","1111110100001011","1111110100111011","0000000010010100","0000001000101001","1111111101110011","1111110111110010","0000000010110011","0000001000011100","1111111110001001","1111111000110110","1111111111100001","0000000001100111","1111111101110010","1111111111000100","0000000000111111","1111111101110100","1111111101110011","0000000010110001","0000000101001100","0000000110100111","0000001000101100","0000000011100011","1111111010100100","1111111011110100","0000000010110000","0000000000010011","1111111001000100","1111111000100111","1111111010101110","1111111010110001","1111111110011100","0000000100011101","0000000100010001","1111111111011101","1111111101111111","0000000001110100","0000000111100101","0000001001000010","0000000010100110","1111111101011010","0000000010100001","0000000111110101","0000000011001011","1111111111001001","0000000011011100","0000000101101000","0000000011011001","0000000110000100","0000001000001011","0000000000011011","1111111010011111","0000000000110110","0000000111011110","0000000101010110","0000000010001000","0000000001000101","1111111111001110","0000000001101011","0000001010010010","0000001101100000","0000000100111100","1111111010000011","1111110111100010","1111111101010001","0000000010101001","0000000001101000","1111111111010000","0000000001100110","0000000011000000","1111111110111110","1111111101101011","0000000010000000","0000000011000000","1111111111110101","1111111111000001","1111111110010011","1111111100101001","0000000000110100","0000000110000111","0000000001010101","1111111001100111","1111111010001110","1111111100100010","1111111011001110","1111111101101111","0000000010111011","0000000100001000","0000000110111011","0000001100110010","0000001001110010","1111111111100010","1111111101011110","0000000010100100","0000000011001111","0000000000110001","1111111111110111","1111111110100100","1111111110101000","0000000000110000","1111111110001001","1111111001001101","1111111101011011","0000000110111111","0000001000100110","0000000011101100","0000000000101111","0000000000100001","0000000011001011","0000000111100011","0000000101110011","1111111110011010","1111111101110000","0000000011110011","0000000100000011","1111111111011000","1111111111000000","1111111110111101","1111111000100100","1111110011010000","1111110111000001","1111111110100111","0000000001010000","1111111101111101","1111111010100001","1111111101010010","0000000101100111","0000001010100001","0000000110000010","1111111101111001","1111111010010110","1111111010011111","1111111001000111","1111111000011111","1111111110001001","0000000101100000","0000000101010101","0000000000011011","0000000000000011","0000000001111111","1111111111101111","1111111101000011","1111111101110001","1111111100001110","1111110111101110","1111111001001010","0000000000110100","0000000100101101","0000000010101010","0000000001010001","0000000010010001","0000000010101000","0000000010010010","0000000010100110","0000000010100001","0000000001000001","0000000000010001","0000000010100101","0000000100111011","0000000001111101","1111111100000000","1111111011011111","0000000000100110","0000000010100110","0000000000000011","0000000001010000","0000000111010101","0000001000111001","0000000011100001","0000000000110101","0000000101000011","0000000111100010","0000000011101011","0000000000110110","0000000010010001","0000000000100101","1111111010011110","1111111000101110","1111111101101010","0000000010001101","0000000011010010","0000000011010000","0000000010111101","0000000001100100","1111111101111010","1111111000010101","1111110110000011","1111111001101010","1111111011101010","1111111000011011","1111111001010000","0000000000011101","0000000001101101","1111111010011100","1111110111011110","1111111100001101","1111111111000011","1111111101010101","1111111101011111","0000000001110001","0000000101101011","0000000100110101","0000000001000010","0000000000111100","0000000101101001","0000000111110000","0000000011111101","1111111111011010","1111111110001001","1111111111111101","0000000011101111","0000000110100001","0000000110011000","0000000100101111","0000000000101111","1111111010101011","1111111010110001","0000000001000001","1111111110110110","1111110101000111","1111110111010001","0000000010010110","0000000000111101","1111111001101000","0000000001001000","0000001101000110","0000001001111010","0000000000110110","0000000000010010","0000000011000000","0000000011001000","0000000010010000","1111111111101110","1111111101110111","1111111110111010","1111111011010011","1111110101000011","1111111100000110","0000001001100011","0000000101000111","1111110111110110","1111111100100011","0000001001100110","0000001000110100","0000000100000001","0000000110011011","0000000100111000","0000000000101001","0000000110011001","0000001010010001","1111111111011011","1111110111110010","1111111110011100","0000000010101010","0000000000100000","0000000100001101","0000000110001110","1111111101001010","1111111001010110","0000000001110011","0000000011011001","1111111011101101","1111111101011110","0000000101111100","0000000100010001","1111111100010111","1111111001101101","1111111011011011","0000000000100110","0000000111001111","0000000011110010","1111111000010100","1111111001001111","0000000111100000","0000001110000010","0000001001010101","0000000101111000","0000000011100011","1111111111010010","0000000000100000","0000000111001011","0000001001111000","0000000111110111","0000000100001110","1111111110100001","1111111100000111","1111111111101110","1111111111100110","1111111100011110","0000000011110011","0000001100011000","0000000010011100","1111110101010111","1111111101011011","0000001010011011","0000000110100011","0000000001011010","0000001000011001","0000001001100101","1111111101101000","1111110111101001","1111111101110001","0000000001000101","1111111011100101","1111110110001100","1111111000010010","1111111111000011","0000000001000110","1111111100001101","1111111001011110","1111111011000111","1111111001000110","1111110111100011","0000000000010000","0000000111111001","0000000000010010","1111110110101000","1111111010100010","0000000010001111","0000000010101110","0000000000111110","1111111111101101","1111111101101110","1111111111101101","0000000011111111","0000000001110000","1111111101101101","0000000001011101","0000000101011010","0000000001011010","1111111110010111","0000000001011001","0000000011001000","0000000011001101","0000000101011010","0000000100010110","1111111111100000","0000000000001000","0000000011011101","1111111111111101","1111111100101101","0000000001110100","0000000011100010","1111111100000010","1111111001111111","0000000001010111","0000000100110000","0000000011010111","0000000100110111","0000000011001101","1111111011110000","1111111011110100","0000000011101101","0000000011000110","1111111011111111","1111111100100001","1111111110010111","1111111000001100","1111110111000101","0000000001101011","0000000110001111","1111111110010000","1111111010000000","1111111110011001","1111111111110011","1111111100101110","1111111100100010","1111111111011010","0000000010000101","0000000010000011","1111111100100001","1111110111010111","1111111100111011","0000000110100011","0000000100111101","1111111101000110","1111111101101001","0000000010100000","0000000001000000","1111111101100100","1111111110100101","1111111111101100","1111111111010100","0000000001001001","0000000011010000","0000000010101110","0000000010001101","0000000001100111","1111111110000111","1111111010111111","1111111010110001","1111111001111100","1111111011010110","0000000101000101","0000001110011010","0000001011011000","0000000011101011","0000000011011010","0000000101010001","0000000001001000","1111111100000001","1111111011101010","1111111110100110","0000000010011110","0000000100001001","0000000001100011","1111111111011011","1111111111110010","1111111011110011","1111110100110000","1111110110011100","0000000000011010","0000000110001111","0000000101011101","0000000011100011","0000000001101100","0000000001010011","0000000011000001","0000000000100001","1111111010000111","1111111010010101","1111111110001100","1111111000111101","1111110010100110","1111111010100001","0000000101010000","0000000001011011","1111111010111101","0000000010001110","0000001011100000","0000000111000101","1111111101100101","1111111100110100","0000000001011001","0000000010110011","0000000001111111","0000000010011100","0000000010010101","1111111111100110","1111111101000010","1111111110100001","0000000011010111","0000000101110000","0000000010001010","1111111110000010","1111111111111001","0000000010110101","1111111111011000","1111111011101111","1111111111110011","0000000011001101","1111111110010101","1111111010110011","1111111101011001","1111111100100001","1111111001011001","1111111111000111","0000000110010010","0000000001011111","1111111010001010","1111111101011000","0000000010101010","0000000000011010","1111111011111000","1111111000100111","1111110101010100","1111110110001110","1111111100001111","1111111111101100","1111111110110001","1111111111001110","0000000000111101","1111111111011110","1111111100000111","1111111100011100","0000000010011110","0000001001010000","0000001001110000","0000000101100001","0000000011100011","0000000010001010","1111111101001101","1111111011111000","0000000010010011","0000000100110111","1111111101111101","1111111001101001","1111111110011011","0000000100001001","0000000100010101","1111111111111001","1111111011011100","1111111101110101","0000000100110001","0000000100100000","1111111111001100","0000000010101000","0000001001100010","0000000101001001","1111111110010011","0000000010100010","0000000101000110","1111111011101111","1111110111100001","0000000001000001","0000000101011100","1111111101001100","1111111010000000","0000000010100101","0000000111001000","1111111111111110","1111111001101110","1111111110100100","0000000110100111","0000000101110010","1111111111110001","0000000000111110","0000000111101001","0000000110111110","1111111111110100","1111111101010000","1111111101011010","1111111000100010","1111110101010000","1111111010111000","0000000000010001","1111111110100000","1111111110010000","0000000010111101","0000000011011100","1111111110011010","1111111101000101","0000000000111001","0000000011101110","0000000011101011","0000000010001110","0000000000111011","0000000001101110","0000000010001110","1111111110001101","1111111001101100","1111111010111000","1111111110000111","1111111110110000","1111111111110100","0000000001111010","0000000010000100","0000000010111101","0000000100101010","0000000000101000","1111111011101110","0000000010001010","0000001100010011","0000001010111100","0000000101101110","0000000111100101","0000000110000011","1111111100010000","1111111001011111","1111111111110100","0000000000101001","1111111101100001","1111111111111101","0000000000101001","1111111100000001","1111111110101010","0000000110010011","0000000010110111","1111111010101011","1111111100111001","0000000000010011","1111111011100100","1111111100011011","0000000101100010","0000000100110010","1111111011110111","1111111101111110","0000000111001100","0000001000000000","0000000101000000","0000000101010010","0000000010110000","1111111111110001","0000000100001010","0000000110010010","1111111110011011","1111111010111011","0000000010010110","0000000101101000","0000000000011100","1111111101111000","1111111101010001","1111111000110011","1111110111101100","1111111101101111","0000000001110100","0000000001010001","0000000001001001","1111111111010100","1111111010010010","1111111001110110","0000000000001010","0000000100101111","0000000011100001","0000000001010101","0000000010001100","0000000100001001","0000000001101100","1111111010100011","1111110111011001","1111111011101111","1111111110010000","1111111010111010","1111111010110110","0000000000101101","0000000011010101","1111111111111001","1111111100111110","1111111110010011","0000000001111111","0000000011101110","0000000001010001","0000000000001011","0000000100001100","0000000100010011","1111111100101001","1111111010111110","0000000010111111","0000000011001101","1111111000110001","1111110111110001","0000000011111010","0000001001110101","0000000010100110","1111111010111001","1111111011000110","1111111111110001","0000000010000111","1111111111101110","1111111110011011","0000000010011001","0000000011111110","1111111110110100","1111111101100001","0000000011101010","0000000100000110","1111111100000100","1111111001000110","1111111100111100","1111111100111101","1111111011100000","0000000001000000","0000000110011111","0000000001111111","1111111010000000","1111111001001101","1111111110010011","0000000010111101","0000000101000110","0000000011111010","1111111111000010","1111111010000000","1111111000111000","1111111011010010","1111111110101111","0000000001001110","0000000000100010","1111111110010101","0000000001001010","0000001000011011","0000001000110010","0000000000110011","1111111111010111","0000000111000001","0000000110010011","1111111010111010","1111111000110111","0000000010011111","0000000011000111","1111111000110000","1111110110111011","1111111111001110","0000000001000101","1111111010111101","1111111001001100","1111111110110100","0000000110000000","0000001001111100","0000000111000010","1111111111001100","1111111010110010","1111111011110001","1111111100001000","1111111100001011","1111111111111101","0000000010111111","0000000001001101","0000000000100100","0000000010101010","0000000000100010","1111111100101101","1111111111110101","0000000011000111","1111111011101001","1111110010111100","1111110110101100","1111111110111100","1111111110010010","1111111001110101","1111111100101110","0000000100110101","0000001001010110","0000000111100010","0000000011010100","0000000010001101","0000000100110111","0000000110001101","0000000011111100","0000000001100100","0000000000110111","0000000000111001","0000000001101100","0000000001001100","1111111101110011","1111111101111111","0000000101100110","0000001001111101","0000000100100010","0000000000110101","0000000100001011","0000000001100010","1111110110111100","1111110110001010","0000000010000111","0000000111000001","1111111110010001","1111111000100010","1111111110000010","0000000010111000","1111111111101101","1111111100111010","0000000000110010","0000000101111011","0000000110111000","0000000100010010","1111111111110001","1111111100100111","0000000000000000","0000000110100100","0000000110010011","0000000000100011","1111111111111111","0000000011101001","0000000010111110","0000000000111011","0000000011011111","0000000100110111","0000000000111001","1111111110011001","1111111111100010","1111111111010000","1111111111010111","0000000010011101","0000000001010111","1111111010010011","1111111001001001","0000000001010001","0000000101111111","0000000010001001","1111111111000110","0000000000110010","0000000001010101","1111111111011100","1111111111111001","0000000011101110","0000000111111111","0000001010100000","0000001001110100","0000000101101101","0000000001101010","0000000001010101","0000000011010011","0000000010110000","1111111110000100","1111111001101110","1111111010101101","1111111110011101","1111111110010101","1111111010100101","1111111001010000","1111111011101110","1111111110110100","0000000001000000","0000000001110001","0000000010011000","0000000110010111","0000001001101101","0000000010111001","1111111000011110","1111111011011100","0000000110111101","0000000111010101","1111111110111100","1111111110000111","0000000010111111","0000000011000000","1111111111001001","1111111010010001","1111110101110110","1111111000111111","0000000001100100","0000000001101001","1111111100101101","0000000010111100","0000001100110000","0000000111101100","1111111011101111","1111111000111011","1111111010011100","1111111010000110","1111111101010111","0000000001100011","1111111111000111","1111111101000101","0000000010000111","0000000011110101","1111111100100001","1111111000111000","0000000000000101","0000000101101101","1111111111101011","1111110111111010","1111111011100110","0000000101001010","0000000110010000","0000000000000001","1111111101110110","1111111111001110","1111111100111101","1111111010000100","1111111100000000","1111111111101000","0000000001101001","0000000010011010","0000000000101010","1111111110110110","0000000001111100","0000000011110101","1111111100110001","1111110111010000","1111111110001111","0000000101110101","0000000010011010","1111111111000110","0000000101001100","0000001001001110","0000000010101101","1111111011111011","1111111110101101","0000000110001111","0000001001110111","0000001000100101","0000000110101100","0000000110110100","0000000111010100","0000000101101011","0000000010000110","1111111111001011","1111111110111111","0000000000001101","1111111111101000","1111111101111100","1111111110000111","1111111101100011","1111111010111011","1111111110110010","0000001010011100","0000001101010011","0000000010101001","1111111110010001","0000000101010011","0000000011000010","1111110101110001","1111110100001001","1111111110010111","1111111111010111","1111110111101101","1111110111010101","1111111101011101","0000000001101111","0000000100010001","0000000011100011","1111111110010010","1111111011111100","1111111110101110","1111111111001100","1111111110111000","0000000011101101","0000000110011100","0000000001111001","0000000000000001","0000000100001001","0000000101000100","0000000010010011","0000000001001010","1111111111000110","1111111101001101","0000000001000001","0000000010100101","1111111011000010","1111111001100000","0000000110100011","0000001110110110","0000000111110100","0000000001111100","0000000100100011","0000000011100110","1111111110010001","1111111101110010","1111111110101101","1111111100100000","1111111110110110","0000000110011010","0000001000001111","0000000100101101","0000000101010011","0000000110110011","0000000000111100","1111111001001101","1111111000110100","1111111101111110","0000000011000111","0000000110010001","0000000101100001","0000000000110000","1111111100010010","1111111011000111","1111111100111011","0000000001101001","0000000110010111","0000000100110101","1111111110001001","1111111011110110","0000000000011011","0000000011000011","1111111111011010","1111111100110010","0000000000101110","0000000100100111","0000000000001100","1111111000001001","1111110111100101","1111111110100000","0000000011000000","0000000001111111","0000000000111000","0000000001110111","0000000001111010","0000000000000011","1111111110011001","1111111111100110","0000000100001000","0000000111110100","0000000110010001","0000000001010111","1111111101010011","1111111011000110","1111111011100111","1111111110101000","1111111111001010","1111111011101001","1111111010101001","1111111110010111","0000000000011000","1111111110101111","1111111101010010","1111111100000001","1111111001101101","1111111000111111","1111111011011100","1111111111010100","0000000001110010","1111111111111110","1111111100110001","1111111110101011","0000000000111010","1111111010010100","1111110100010010","1111111011010001","0000000011010010","1111111111111110","1111111110000001","0000000011011100","0000000000010100","1111110101100100","1111110111011011","0000000010010100","0000000010010100","1111111011101011","1111111100111000","0000000000000101","1111111101111000","1111111111001010","0000000110100000","0000001000000011","0000000001001001","1111111100010010","1111111100110110","1111111101000000","1111111101010100","0000000010110111","0000000111111111","0000000010101000","1111111001000100","1111111010010111","0000000011000110","0000000100010001","1111111111111110","0000000001001000","0000000010011001","1111111011100000","1111110110010010","1111111100011110","0000000101000001","0000000101101000","0000000010000000","0000000001010100","0000000100011101","0000000111011101","0000000101100100","1111111111111100","1111111110010000","0000000010000011","0000000011011010","1111111111111010","1111111110101000","0000000001001010","0000000000010101","1111111011000100","1111111010000010","1111111111100011","0000000001101001","1111111011010111","1111110110010101","1111111001110011","1111111110111111","0000000000010100","0000000010010000","0000000101000111","0000000010011110","1111111100100110","1111111011110101","1111111111101011","0000000010111010","0000000101010010","0000000101110000","0000000001000111","1111111011101111","1111111100110100","0000000001001110","0000000001000010","1111111101110011","1111111110001000","0000000000101110","1111111111001000","1111111010100101","1111111011010001","0000000001001001","0000000001111011","1111111011101010","1111111001000010","1111111101010000","0000000000001011","0000000001010001","0000000101110101","0000000110110001","1111111101000010","1111110110010001","1111111111001110","0000001001110111","0000000101001010","1111111010110010","1111111100001100","0000000110000011","0000001001101110","0000000011110011","1111111100011000","1111111001110000","1111111010001001","1111111001000010","1111110111010111","1111111000101101","1111111011101011","1111111101110001","0000000000100010","0000000010111001","0000000000101100","1111111101100101","1111111111111101","0000000010111011","0000000000000101","1111111101011001","1111111111011101","1111111111111101","1111111100110011","1111111011001000","1111111011001001","1111111100101100","0000000010111100","0000000110100011","1111111110000001","1111110101001001","1111111010100001","0000000001110110","1111111100111100","1111111000110110","0000000001101100","0000001010001101","0000000111010000","0000000010011000","0000000011001010","0000000011101101","0000000000010110","1111111110000001","1111111110110100","1111111101010111","1111110111001101","1111110100011100","1111111010011110","1111111111010011","1111111011100101","1111111010110110","0000000011100110","0000000111010110","0000000000110100","1111111111110001","0000000111100101","0000001001011110","0000000011101110","0000000000011001","1111111110101010","1111111011111101","1111111110011111","0000000101001100","0000000110111001","0000000011010001","1111111111010100","1111111101001100","0000000001101110","0000001100100010","0000001111110001","0000000110010111","1111111110110001","1111111111001110","1111111110101000","1111111110010110","0000000110011001","0000001101101101","0000001000010111","1111111110010100","1111111100000001","0000000000001111","0000000011111101","0000000010101010","1111111100001011","1111111000010101","1111111101011001","0000000011010111","0000000001000110","1111111100000010","1111111011101111","1111111101110110","0000000000001111","0000000100011001","0000000110101011","0000000011011111","0000000000100100","0000000011001000","0000000101100101","0000000001101010","1111111011111011","1111111101011100","0000000110010010","0000001100111010","0000001011000110","0000000101010010","0000000001001010","1111111101110101","1111111011000100","1111111100101001","0000000001000000","0000000001000000","1111111101100011","1111111111110001","0000000111110011","0000001001010011","1111111111010000","1111110110111011","1111111011011000","0000000010010011","1111111110100101","1111111001000011","1111111110111010","0000000111110101","0000001000000000","0000000110011011","0000001001011110","0000001000101001","0000000010000011","1111111111101000","0000000001000011","1111111110101001","1111111100110010","0000000001001010","0000000011001100","1111111011110001","1111110011010101","1111110100011110","1111111110001000","0000000110111011","0000000111100101","0000000010001100","1111111101110101","1111111011101001","1111111001101001","1111111011010010","0000000001000111","0000000011101011","0000000010001010","0000000100101010","0000001001011100","0000000111001011","0000000000111010","0000000000011110","0000000011010001","0000000000111011","1111111011100011","1111111011010101","0000000001011101","0000000110111110","0000000100101111","1111111100100111","1111111000110111","1111111101101100","0000000001110110","1111111110011100","1111111100000010","0000000011000000","0000001010010000","0000000110010111","1111111101110011","1111111011100101","1111111011111110","1111111001101100","1111111010110100","1111111111010101","1111111101101001","1111111010011100","0000000001000010","0000000110111101","1111111110110110","1111110110100101","1111111011110101","0000000001011001","1111111110011011","1111111110101111","0000000011111101","0000000011001011","1111111111110101","0000000001101000","0000000010001011","1111111111011100","0000000010010011","0000001000000100","0000000110010111","0000000000101000","1111111111000010","1111111111010011","1111111110010110","1111111110100100","0000000000000000","0000000000001101","1111111101101110","1111111000101110","1111110110001010","1111111010111111","0000000001010001","0000000001000001","1111111101001100","1111111001100100","1111110101010011","1111110110110010","0000000010100110","0000001010011011","0000000010111000","1111111001101001","1111111011000000","1111111100101000","1111110110110010","1111110010110010","1111110110000011","1111111010111110","1111111110110110","0000000010011011","0000000100001111","0000000100101111","0000000101101000","0000000100011111","0000000001010000","0000000001110110","0000000111000000","0000001010000111","0000001001001111","0000000111001011","0000000011010010","1111111111100000","0000000010100100","0000001000110101","0000000101001110","1111111001100100","1111110110101110","1111111111001110","0000000100011111","0000000000110111","1111111100011000","1111111100001100","1111111110010100","1111111110110011","1111111011010110","1111111000111100","1111111110000101","0000000100000011","0000000001101000","1111111110011011","0000000010111101","0000000110110100","0000000101110000","0000001000100110","0000001011111011","0000000100001011","1111111010010001","1111111100100100","0000000011010110","0000000011100111","0000000010010101","0000000100011000","0000000111010111","0000001001101001","0000000110010110","1111111011110000","1111110111001100","1111111110001110","0000000000000000","1111111001101011","1111111111010101","0000001101011001","0000001010000110","1111111010010101","1111110111111010","1111111111010001","1111111101110100","1111111000011000","1111111001111000","1111111101000101","1111111110101011","0000000011101111","0000000111111100","0000000011001001","1111111011101111","1111111100001111","0000000000110111","0000000000010011","1111111100011010","1111111100010010","1111111110010101","1111111101111011","1111111111000010","0000000101010011","0000001000101100","0000000010111000","1111111011110101","1111111011100100","1111111111011000","0000000010111110","0000000011111001","1111111111111100","1111111100010111","1111111111100111","0000000001110010","1111111011101101","1111111001001010","0000000000101001","0000000011011010","1111111101001111","1111111101100011","0000000100011001","0000000010100000","1111111011000100","1111111011010100","1111111110111100","1111111110100101","0000000000001000","0000000100101000","0000000100000101","0000000000111010","0000000010010011","0000000010110101","1111111101110001","1111111100100000","0000000010101000","0000000011010100","1111111010111111","1111111000110101","0000000000111010","0000000010101010","1111111010100000","1111111010100010","0000000101111111","0000001001110000","0000000010011001","0000000000001011","0000000100011110","0000000011010100","1111111111000010","1111111111100010","0000000000100100","0000000000000000","0000000011101100","0000000111101110","0000000011101001","1111111110010101","0000000010010010","0000001001111101","0000001010001110","0000000011100010","1111111110111101","0000000000010110","0000000000001101","1111111001011011","1111110110111110","0000000000001101","0000000101101101","1111111101011111","1111110111011001","1111111011001001","1111111010110010","1111110110010010","1111111011010000","0000000010101011","0000000000100000","1111111110001111","0000000001001101","1111111111010001","1111111101011100","0000000111001000","0000001110111001","0000001000001101","0000000001100000","0000000010101110","1111111111110000","1111111010011011","1111111110111100","0000000101110001","0000000011111110","0000000001000000","0000000001001101","1111111101111110","1111111010111000","1111111110011100","1111111111110101","1111111001011100","1111110110011001","1111111011010110","1111111110100011","1111111101110101","0000000000010011","0000000100010011","0000000010110111","1111111110111101","0000000000011010","0000000100111100","0000000011100100","1111111100101001","1111111010110010","0000000001011000","0000000111010100","0000000110111101","0000000011110100","1111111110110000","1111110111101000","1111110101111101","1111111100110110","0000000010010001","0000000000100111","1111111110100010","1111111110011011","1111111100110101","1111111100010000","1111111110011101","1111111110100000","1111111100101111","1111111101001011","1111111100000000","1111111000101000","1111111100000011","0000000100101101","0000000110011011","0000000010011100","0000000001001100","1111111111111100","1111111101101000","0000000000110111","0000000100000100","1111111110010110","1111111001110011","1111111101111100","1111111110000111","1111111000001110","1111111011011101","0000000100001001","0000000010010111","1111111101110111","0000000011100111","0000000111010101","1111111110010101","1111110101101001","1111110110100101","1111111010001101","1111111100101110","1111111110001100","1111111010101000","1111110101100011","1111111000001110","1111111111000001","0000000000001001","1111111110001000","1111111110000001","1111111100001011","1111111000110010","1111111001111011","1111111101100000","1111111110010100","1111111111110011","0000000011000101","0000000000001001","1111111000011010","1111111000110101","0000000000101001","0000000001100001","1111111011111100","1111111101000101","0000000010110000","0000000000110100","1111111011010111","1111111101111101","0000000011100100","0000000001011111","1111111100111010","1111111111010010","0000000011110010","0000000010001111","1111111110101001","0000000001000010","0000000111000111","0000001000001101","0000000010100110","1111111101100101","1111111110001000","0000000000111011","0000000010011111","0000000100001110","0000000110011011","0000000110101101","0000000101111000","0000000101111000","0000000100110000","0000000010010000","0000000001111100","0000000010101111","0000000000101101","1111111110010011","1111111110111101","1111111110110111","1111111100000011","1111111011001111","1111111101100010","1111111110110100","1111111111000000","1111111111100000","1111111110111111","1111111111011110","0000000010110110","0000000011010000","1111111111010110","0000000001101011","0000001010111001","0000001011110110","0000000010101010","1111111110010110","0000000000001000","1111111100101110","1111110111111010","1111111100011011","0000000101000010","0000000111001011","0000000011000100","1111111100110101","1111111000110111","1111111100010010","0000000001111001","1111111111000100","1111111001100001","1111111100110111","0000000001110010","1111111111000000","1111111101110011","0000000001101111","1111111101010000","1111110010100101","1111110101010010","0000000011001111","0000000111101111","0000000001001110","1111111101001011","1111111101010011","1111111110001001","0000000010111001","0000001000100001","0000000101111111","1111111111010100","1111111111110011","0000000100010010","0000000011000101","0000000000011100","0000000100010101","0000001000110100","0000000110100101","0000000011111010","0000000101111111","0000000100111011","1111111101101101","1111111010001000","1111111100110110","1111111110000111","1111111110001001","0000000001100100","0000000010110001","1111111110110010","1111111110000110","0000000000110000","1111111101110001","1111111001111110","1111111101010100","1111111110101010","1111111011000010","0000000001011000","0000001101110000","0000001000111000","1111111001100111","1111111011010010","0000000110011111","0000000011001101","1111111100000000","0000000010011110","0000000111001000","1111111110000000","1111111010000101","0000000011000100","0000000110001000","1111111111001101","1111111101000010","1111111111110101","1111111111010011","1111111111110001","0000000011011000","0000000010110011","1111111111111001","0000000001100101","0000000010111110","0000000000010110","0000000000010001","0000000001100000","1111111110001111","1111111110111011","0000000111111111","0000001001011000","1111111111000000","1111111101100010","0000000111111110","0000000111100000","1111111001101111","1111110101110000","0000000000101111","0000001001000100","0000000110011110","0000000000001100","1111111101100111","1111111111111101","0000000001110101","1111111110001001","1111111011010000","0000000000010111","0000000100011111","1111111110111100","1111111011001000","0000000010111001","0000001001101111","0000000100001001","1111111011011111","1111111010110111","1111111111001011","0000000010000000","0000000010010111","0000000001101100","0000000001111100","0000000010101011","0000000000111010","1111111111010101","0000000100000011","0000001010110101","0000001001100000","0000000001100111","1111111100000010","1111111010111000","1111111101011101","0000000011010101","0000000101110001","0000000000111001","1111111101111001","0000000001011011","0000000010100101","0000000000001000","0000000010000001","0000000100000110","0000000000010011","0000000000000111","0000000101111100","0000000011000011","1111111000111100","1111111001011000","0000000000100001","1111111110110111","1111111011100101","0000000000010100","0000000001111010","1111111100101100","1111111101001011","0000000000110000","1111111101010101","1111111101010010","0000000111100111","0000001010011100","1111111111010100","1111111010011010","0000000010000100","0000000101010110","0000000000000110","1111111101110000","1111111111001010","1111111101111100","1111111101101011","0000000011101111","0000001001110100","0000000101011110","1111111000110001","1111110011110001","1111111111100010","0000001101101001","0000001100000011","0000000001101101","0000000000011111","0000000101101000","0000000011011010","1111111100010100","1111111011001111","1111111111010110","0000000010011010","0000000011101001","0000000010000110","1111111101000111","1111111011100101","0000000001110101","0000000101111010","1111111111111001","1111111010000100","1111111110011000","0000000011011001","1111111110101101","1111111000101000","1111111100000001","0000000011000001","0000000011011101","1111111111000010","1111111101110000","0000000010010110","0000000111011010","0000000100100100","1111111010100100","1111110101100001","1111111010110111","0000000001000100","0000000001111001","0000000010011000","0000000011100110","0000000001100000","1111111111001010","1111111111110111","1111111111001110","1111111101111000","0000000001111111","0000000110101000","0000000011010010","1111111101001101","1111111010111100","1111110111111101","1111110011101010","1111110100101101","1111111001001000","1111111100001001","0000000001011011","0000000111010011","0000000101000111","0000000000000101","0000000010111101","0000000110010011","0000000000111000","1111111100010001","1111111111000000","0000000000001100","1111111101111111","1111111110110011","1111111111000001","1111111100001010","1111111111010001","0000000110101101","0000000101001100","1111111110001111","1111111110111001","0000000010011111","0000000001000111","0000000010001111","0000000111011101","0000000101011100","1111111101011110","1111111011001101","1111111100010011","1111111001000111","1111110110001111","1111111000110001","1111111100101000","1111111110001011","1111111101001000","1111111011010011","1111111101110111","0000000011000100","0000000000100101","1111111001111000","1111111101110111","0000000110110111","0000000011100011","1111111011110110","0000000000111001","0000001000111111","0000000101010110","1111111111011000","0000000001000010","0000000010100010","1111111111101010","1111111101011000","1111111010011111","1111110101110101","1111110101101011","1111111010001111","1111111101101110","0000000010100011","0000001010001110","0000001010000110","1111111111000110","1111110111111000","1111111011001010","1111111101011010","1111111010001010","1111111011110000","0000000100011100","0000001001111000","0000001000100100","0000000110010101","0000000100011001","0000000000011010","1111111100101100","1111111100000010","1111111110000101","0000000011000111","0000001000111111","0000001000001100","1111111111010101","1111110111100110","1111110110011100","1111111001000111","1111111110111011","0000000110101010","0000001000001111","0000000001011111","1111111100100101","1111111110111011","0000000001101101","0000000000101100","1111111111010011","1111111110101000","1111111100001011","1111111001010111","1111111010110000","1111111111010001","1111111111100110","1111111011001011","1111111011011000","0000000001011000","0000000001110101","1111111100111010","1111111110111000","0000000010111100","1111111100100000","1111110110111110","1111111111010110","0000000101101111","1111111111101101","1111111111100100","0000001001001011","0000000110101111","1111111001011110","1111111000001010","0000000000111111","0000000011000101","0000000000100111","0000000000101010","1111111111000010","1111111100001000","1111111100100111","1111111100100100","1111111010011011","1111111011101110","1111111110011101","1111111101001001","1111111010110001","1111111001110001","1111111001101000","1111111110101110","0000000111010110","0000001000011110","0000000100001010","0000000100001111","0000000001010011","1111110110001101","1111110100110010","0000000000111000","0000000010101010","1111111000010010","1111111010001101","0000000101100110","0000000011101011","1111111011000110","1111111110011110","0000000100110100","0000000001011011","1111111101110011","0000000001000000","0000000011001001","0000000001010101","1111111111110110","1111111110101010","1111111100111101","1111111100110001","1111111111000011","0000000011101011","0000000101111000","1111111101101110","1111110010101101","1111110110111010","0000000100100111","0000000101000110","1111111100001011","1111111101110110","0000000100000011","1111111111001111","1111111000010111","1111111001110111","1111111010001110","1111110110111111","1111111010010001","1111111111011110","1111111100000100","1111111000011100","1111111110011001","0000000101011101","0000000101011110","0000000010110100","0000000001010111","0000000001000101","0000000010100110","0000000100001111","0000000100011001","0000000101001110","0000000101101110","0000000011111001","0000000100100011","0000000111010010","0000000001100111","1111110110011010","1111110101111100","1111111101110110","1111111101100001","1111110110111011","1111110110100001","1111111010000101","1111111100000110","1111111111101101","0000000011101111","0000000100001101","0000000100000011","0000000010110011","1111111101011100","1111111100111110","0000000101001001","0000000101001001","1111111001101111","1111111001001001","0000000100110101","0000000100010111","1111111001000011","1111111010111001","0000000110100101","0000000110111100","1111111110100010","1111111100001011","1111111111000001","0000000000100000","0000000000110011","0000000000011000","0000000000010100","0000000011011110","0000000110100000","0000000100100010","0000000010001100","0000000011110101","0000000011100001","1111111110001010","1111111011001011","1111111101110010","1111111111100110","1111111110010000","1111111110100111","0000000000110110","1111111111101010","1111111100011110","1111111101110100","0000000010001010","0000000010011101","1111111111100011","1111111110100100","1111111101101000","1111111010000000","1111111000100111","1111111100111101","0000000010000110","0000000011001101","0000000001100101","0000000001001110","0000000011111010","0000000101101100","0000000010000100","1111111110001001","0000000000100101","0000000010111010","1111111111010010","1111111111010001","0000000101100100","0000000011010101","1111111000101000","1111111000100110","0000000001010110","1111111110010111","1111110011100001","1111110100111001","1111111111000101","0000000011001100","0000000100001000","0000000111000100","0000000100001001","1111111100000111","1111111100001110","0000000011110110","0000000101110011","0000000010001101","0000000010001011","0000000011101010","0000000001110111","0000000001100001","0000000011011011","1111111111111110","1111111010011000","1111111101101000","0000000011111111","1111111111111001","1111110111100000","1111111000001000","1111111101001101","1111111110100010","0000000000111001","0000000101000110","0000000011101100","0000000000111011","0000000110100101","0000001101111000","0000001011100100","0000000011111110","1111111111111001","1111111111011100","1111111111010011","1111111100011000","1111110110101010","1111110101111001","1111111101001110","0000000010000001","1111111111101101","1111111111101111","0000000010010011","1111111101101011","1111110110010101","1111110111011001","1111111110000011","0000000100010101","0000001001010000","0000000110011011","1111111100001111","1111111100000000","0000001000011101","0000001011011100","0000000000011000","1111111011101111","0000000000100111","0000000000000000","1111111011110000","1111111110111011","0000000101101100","0000001000101011","0000001000011000","0000000101001100","0000000001010000","0000000001100100","0000000010001001","1111111110000110","1111111101110111","0000000100001010","0000000011010101","1111111010011110","1111111010101010","0000000011110101","0000000100110001","1111111101000100","1111111001101011","1111111100011110","0000000001010100","0000000110010011","0000000100111101","1111111011011101","1111110110010010","1111111011001000","1111111101110100","1111111001110010","1111111001001010","1111111100110001","1111111100000010","1111111001100010","1111111011011001","1111111101001010","1111111100010111","1111111110001110","0000000001000001","1111111111100011","1111111110100011","0000000001010100","0000000001011010","1111111111010111","0000000001111110","0000000011110000","1111111110010100","1111111011010000","1111111110101010","1111111100111110","1111110111111100","1111111101010111","0000000100111010","1111111110010000","1111110110000000","1111111101100101","0000000110111001","0000000000111011","1111110110111111","1111110111010101","1111111100110011","0000000000000011","0000000000101110","1111111101000010","1111110111100000","1111111010011000","0000000101011100","0000001010110100","0000000110111010","0000000101100100","0000001001000001","0000000101101001","1111111100010101","1111111100001010","0000000100011011","0000000100111001","1111111110000001","1111111101000011","1111111110111111","1111111011111001","1111111101000111","0000000110010101","0000000111011000","1111111110010001","1111111101101011","0000000101010010","0000000011101111","1111111100111101","1111111111010110","0000000011101110","1111111110101101","1111111000000100","1111111000001010","1111111010011111","1111111100101110","0000000001010010","0000000011101010","1111111110001111","1111110111000001","1111111000101011","0000000001111010","0000000101100001","1111111101111001","1111110110101110","1111111010000011","0000000000010111","0000000000000100","1111111100110100","1111111101011101","0000000010010101","0000000111110101","0000001000101110","0000000100001011","0000000000111101","1111111111001010","1111110111101011","1111110011010101","1111111111100010","0000001100001111","0000000101010001","1111111011111100","0000000010101001","0000000101111111","1111111010011101","1111110110110100","0000000000011100","0000000001110111","1111111100111000","0000000001010010","0000000100100111","1111111100110100","1111111010110010","0000000011111100","0000000110011111","0000000001000010","0000000000111001","0000000011010100","0000000010101110","0000000101010100","0000001000010101","0000000010011101","1111111100110011","0000000010011001","0000000111101000","0000000001011001","1111111010110001","1111111110110011","0000000110010111","0000000110010111","1111111110111010","1111111001100111","1111111101000111","0000000010110100","0000000001001110","1111111101011011","0000000000111000","0000000111001001","0000001000000111","0000000101111011","0000000100001011","0000000011011100","0000000110001011","0000001001011101","0000000101001010","1111111101111101","1111111111100111","0000000101100101","0000000101010011","0000000011110101","0000000110100110","0000000101010110","1111111111000100","1111111110000110","1111111111111010","1111111010101111","1111110101111101","1111111100000101","0000000011001111","0000000000011111","1111111100101000","0000000000111111","0000000110100001","0000000110101000","0000000110100101","0000001001000100","0000000111100101","0000000000100001","1111111100110010","0000000001011110","0000000110111011","0000000100101101","1111111110100100","1111111110000000","0000000010111100","0000000100010010","1111111110111010","1111111010100101","1111111100101100","0000000000011000","0000000000110100","0000000000101100","0000000001000000","1111111110001101","1111111010101011","1111111011110001","1111111101110010","1111111100001111","1111111100101010","1111111111110101","1111111100001000","1111110100100111","1111110111101000","0000000000101010","0000000000100010","1111111101010001","0000000010100101","0000000110000111","1111111111101000","1111111100111111","0000000011011001","0000000100000011","1111111101010110","1111111101010111","0000000011000111","0000000010111100","1111111111011101","0000000000011101","0000000010010111","0000000001011100","0000000001000011","1111111111111101","1111111010010001","1111110110001100","1111111011111001","0000000100100100","0000000100001101","1111111110110111","1111111111110101","0000000011010000","1111111111110101","1111111100111001","0000000010100110","0000000100101101","1111111011100000","1111110111110100","0000000000101110","0000000011011111","1111111011111010","1111111100011111","0000000011100111","1111111111100100","1111111000011001","1111111111001111","0000001000000001","0000000011001001","1111111101000010","0000000010001010","0000000111111111","0000000100111101","1111111110110100","1111111100101101","0000000000100100","0000000110111011","0000000111001010","0000000000110111","1111111111010000","0000000011110010","0000000011000001","1111111100101101","1111111010111100","1111111101001000","1111111101110000","0000000000110011","0000001000000100","0000001011000101","0000000111010101","0000000101000101","0000000110111100","0000000101100000","1111111101110110","1111111000101111","1111111101101010","0000000100101011","0000000010001101","1111111100110111","0000000001001101","0000000110110001","0000000000100010","1111111001110110","1111111110111111","0000000011011100","1111111111110000","0000000001010101","0000000111101011","0000000011101101","1111111101011011","0000000011011101","0000000110101001","1111111010110000","1111110101000100","1111111111011010","0000000010100101","1111111001011011","1111111011001000","0000001000000011","0000001001010011","1111111111111110","0000000000001111","0000001010001110","0000001101111000","0000001000010111","0000000100111110","0000001000010011","0000001001011101","0000000001110111","1111111001110001","1111111001111000","1111111100101110","1111111101011111","0000000001011101","0000000101010001","1111111111011001","1111111001011110","0000000000111100","0000000111101101","1111111101110010","1111110010111001","1111111000001101","0000000001011111","0000000001000000","1111111110011110","0000000001011011","0000000100101000","0000000011100111","1111111111110000","1111111011111001","1111111011101000","1111111111011000","0000000001101100","1111111111101100","1111111101011101","1111111110100111","0000000001011010","0000000010000011","0000000001011000","0000000101001010","0000001100101110","0000001101111000","0000000111101111","0000000110111000","0000001011100001","0000000111001111","1111111100000111","1111111010111101","0000000010101010","0000000101000010","0000000010011000","0000000001100110","1111111111010111","1111111010100100","1111111010111001","0000000000111110","0000000101000001","0000000100100011","0000000001011110","1111111011111111","1111110110111000","1111110111000000","1111111010101010","1111111011010101","1111111000000001","1111110110101110","1111111100011010","0000000110011111","0000001100010110","0000000111101100","1111111100011001","1111110110100100","1111111100001111","0000000011100111","0000000001100101","1111111100110010","0000000000101001","0000000110000110","0000000001001010","1111111001100111","1111111100101001","0000000100001110","0000000100001000","1111111111001010","1111111110000010","1111111111111010","1111111111110011","1111111110011100","1111111111110011","0000000011000100","0000000100010011","0000000100101111","0000000111010101","0000000111100000","0000000010010111","0000000000011100","0000000100001010","0000000010000111","1111111010111001","1111111100110101","0000000011101000","1111111110011111","1111110011100011","1111110011110101","1111111011101001","1111111111110000","0000000000011001","1111111111001000","1111111101000001","1111111110101000","1111111111110110","1111111001111010","1111110111001101","0000000000000001","0000000101101111","0000000000111110","0000000000100010","0000000101100001","0000000001001000","1111111001011010","1111111101000011","0000000011010000","0000000001100101","0000000001100101","0000000101110101","0000000010110110","1111111011111011","1111111101101001","0000000010110110","0000000010000000","0000000001101001","0000000110100100","0000001000000001","0000000010111110","1111111111111101","0000000001010011","0000000000110010","1111111101000110","1111111010110001","1111111100000110","1111111110011100","1111111101011111","1111111010001111","1111111100011101","0000000011111110","0000000011011100","1111111001011101","1111111000001101","0000000010100010","0000000011110011","1111111010100110","1111111100010101","0000000110011010","0000000011101110","1111111011100101","0000000000101010","0000000110101001","1111111111000101","1111111010010010","0000000010010001","0000000110110001","0000000011111010","0000000110011001","0000001001110101","0000000100011010","0000000000001101","0000000011010111","0000000010010001","1111111100011000","1111111110000111","0000000100011010","0000000011110010","1111111111011011","1111111110101100","1111111111110100","0000000000111110","0000000010011011","0000000000110001","1111111100011001","1111111011001101","1111111100110110","1111111100101111","1111111100110110","1111111111111111","0000000010110000","0000000001111111","1111111110101011","1111111011000100","1111111011010101","0000000000101001","0000000010111011","1111111100111111","1111111000110011","1111111110111110","0000000110000100","0000000010110111","1111111010101000","1111110111110010","1111111010011000","1111111100100011","1111111100110011","1111111110010111","0000000010101100","0000000101010001","0000000001111011","1111111101000011","1111111100111010","1111111111001101","0000000000011001","0000000011011101","0000001000000110","0000000111100111","0000000010100000","1111111111101111","1111111101110101","1111111000110001","1111110111011101","1111111110000100","0000000001100001","1111111100010110","1111111010010101","1111111111100000","0000000000001000","1111111100110001","0000000010101101","0000001011110010","0000000110110101","1111111100101101","0000000000000011","0000000110000001","1111111101111011","1111110110100010","1111111111010001","0000001000010001","0000000100111011","0000000001110001","0000000011011100","0000000000110000","1111111110111101","0000000101010100","0000000110100011","1111111100100111","1111111000100100","1111111111010111","0000000001100011","1111111100010100","1111111010010011","1111111100101110","0000000000110011","0000000110011100","0000000111000100","0000000000011100","1111111110110100","0000000101000100","0000000100000010","1111111001100010","1111110101011011","1111111010001101","1111111011001111","1111111000000110","1111111011000110","0000000010010011","0000000010001001","1111111011110101","1111111101011110","0000001000010101","0000001011100110","0000000010110110","1111111110101000","0000000010100101","1111111111011101","1111110110100111","1111110111101011","1111111101101100","1111111011101100","1111111001111001","1111111111101111","0000000001110101","1111111110111001","0000000011010111","0000001010001010","0000000110100000","0000000000000011","0000000000001101","1111111111100110","1111111100010110","1111111110001110","0000000001001011","1111111110010111","1111111101010010","0000000001000111","1111111111001110","1111110111101100","1111110110011000","1111111010000100","1111111001011011","1111111000001110","1111111101100100","0000000100010000","0000000110010011","0000000110001111","0000000101010001","0000000011011001","0000000110001000","0000001100101101","0000001010101110","1111111111001110","1111111010101101","0000000001001100","0000000011101000","1111111110110110","1111111110011110","0000000010011101","0000000011101010","0000000101011111","0000000111111101","0000000010011100","1111111010111111","1111111110111011","0000000110000011","0000000011011111","1111111111111101","0000000010010010","0000000001000110","1111111101111001","0000000001101010","0000000011001001","1111111011111101","1111111011100110","0000000011101000","0000000000100001","1111110110100000","1111111010000010","0000000001010110","1111111010000111","1111110011001000","1111111011001011","0000000000100111","1111111001011110","1111111000110000","0000000011111111","0000000111011010","1111111110111100","1111111101000111","0000000110010101","0000001010000011","0000000010000110","1111111100010101","0000000000111000","0000000100111101","0000000000010101","1111111100001100","0000000000000011","0000000100000001","0000000010000001","1111111111011011","1111111110010110","1111111011100000","1111111001110111","1111111100010101","1111111101110100","1111111101001111","0000000000000000","0000000011001011","1111111111101010","1111111010010101","1111111010111001","1111111101111001","1111111110100111","1111111110101111","1111111110000100","1111111011101010","1111111011110001","1111111111100001","0000000010011100","0000000101000010","0000001000101011","0000000111001011","0000000000100110","1111111111011111","0000000001110100","1111111011010101","1111110011011110","1111111010010111","0000000110001100","0000000101011010","0000000001000101","0000000110001100","0000001001111010","0000000011010101","1111111101010101","1111111101000110","1111111011010011","1111111000101001","1111111010001100","1111111100000011","1111111011110010","1111111100010000","1111111011001111","1111111000111001","1111111101001100","0000000101001011","0000000100011100","1111111110100001","1111111111011010","0000000011000101","0000000001111000","0000000000101110","0000000001010100","1111111110011111","1111111100101010","0000000001010101","0000000101010001","0000000010111110","1111111111100100","1111111110011100","0000000000010111","0000000101111100","0000001000010000","0000000011011011","0000000010001100","0000000110100101","0000000010001011","1111111000100101","1111111100101001","0000000101111001","0000000000011111","1111111000110100","1111111111011010","0000000100000101","1111111011010100","1111110111011111","1111111111111001","0000000100100011","0000000010011011","0000000010010010","0000000000000000","1111111001110001","1111111011110011","0000000100101101","0000000010111111","1111111001001011","1111111011011111","0000000110111011","0000000100010011","1111110100110010","1111110010000000","1111111111110000","0000000110101100","0000000000011100","1111111110101100","0000000011101101","0000000000011110","1111111000011011","1111111010111011","0000000011000110","0000000101001010","0000000101001011","0000000101101001","0000000000100101","1111111100101100","0000000010111000","0000000111010000","0000000000111110","1111111101010101","0000000000010011","1111111100100110","1111110110110000","1111111110001111","0000001000110010","0000000101101001","1111111111110011","0000000100100010","0000001000101001","0000000011001011","1111111110000001","1111111110000110","1111111101101110","1111111110011010","0000000011011010","0000000101010111","0000000000010001","1111111101011000","0000000000101111","0000000000110000","1111111010100101","1111111010000010","0000000011000100","0000001000000000","0000000001110100","1111111100010100","1111111111011010","0000000010111000","0000000010001100","0000000010111000","0000000011110111","1111111111111111","1111111101100110","0000000010100010","0000000101101001","0000000001001000","1111111110100011","0000000001110101","0000000001101001","1111111100010100","1111111010110101","1111111110000010","1111111111100111","0000000000010101","0000000011001010","0000000011000111","1111111101000110","1111111000111010","1111111100011111","0000000001000011","0000000000010000","1111111110110001","1111111111010000","1111111011111000","1111110110100101","1111111010001011","0000000011101101","0000000100100001","1111111101111101","1111111101110101","0000000011000111","0000000010011111","1111111101010110","1111111100100101","1111111111110111","0000000001011100","0000000000001011","1111111111010110","0000000001100010","0000000011111111","0000000001010101","1111111100001001","1111111101000001","0000000011000100","0000000100100000","1111111110110110","1111111001011011","1111111010110110","0000000001111011","0000000101111100","0000000001000100","1111111011011001","1111111110011101","0000000011001001","1111111111100010","1111111010010010","1111111100011101","0000000001101111","0000000100010010","0000000101011100","0000000110100110","0000000111110000","0000000111111100","0000000011000111","1111111010110000","1111111000100110","1111111101011010","1111111111001010","1111111101110110","0000000000010111","0000000010000010","1111111101001110","1111111001100111","1111111011101101","1111111101001100","1111111101011111","0000000000010011","0000000000000100","1111111001110101","1111110111011111","1111111101100111","0000000011101011","0000000100110111","0000000011101000","0000000000100110","1111111110101000","0000000010111011","0000000111101110","0000000010011000","1111111000011010","1111110111000111","1111111100001111","1111111101100101","1111111101000101","0000000001100001","0000000111000011","0000000110110011","0000000010101000","0000000000000001","0000000000100001","0000000011001000","0000000101111001","0000000101111110","0000000011000011","0000000000100111","0000000000100001","1111111111100111","1111111011100101","1111111000001011","1111111001100101","1111111101100110","0000000000111110","0000000101100110","0000001010111000","0000001001111111","0000000010101100","1111111110011111","0000000000010101","0000000001001110","1111111111011100","1111111111101110","0000000001110010","0000000010101010","0000000010111010","0000000010011100","0000000000001000","1111111101100101","1111111011001101","1111111000010100","1111111001001011","1111111110110000","0000000000010101","1111111100110101","1111111111000110","0000000101110000","0000000011001101","1111111010110000","1111111100001101","0000000100101100","0000000101000110","1111111111000100","1111111111000011","0000000100110000","0000000110110100","0000000011111101","0000000001010111","0000000000000101","1111111110101000","1111111111011101","0000000011010011","0000000011001011","1111111100101010","1111111010001010","0000000000010110","0000000100010010","0000000000010000","1111111011101111","1111111001101010","1111111000111110","1111111111001001","0000001000110100","0000000111000110","1111111101000100","1111111100101100","0000000011100010","0000000010111100","1111111110001100","1111111100110111","1111111010111001","1111111010101101","0000000001111111","0000000100101011","1111111011100011","1111111001100010","0000000110000001","0000001010010010","1111111101111011","1111110110100111","1111111110011011","0000000101111111","0000000010101100","1111111010001110","1111110100111110","1111110110000101","1111111011000010","1111111110010010","1111111101010110","1111111010001001","1111111001000010","1111111110111110","0000001000010000","0000001000000111","1111111101111111","1111111001001001","1111111100011111","1111111011011011","1111110111110000","1111111110001010","0000000111110000","0000000101001111","1111111101100001","1111111110111101","0000000100000001","0000000010001111","1111111110110101","0000000001001101","0000000101001111","0000000101100111","0000000011110010","0000000010001010","0000000000111000","1111111111011100","1111111100111000","1111111001110001","1111111001101011","1111111101011110","0000000000100101","0000000000101011","0000000001001010","0000000010110111","0000000001011111","1111111101000001","1111111011111101","0000000000000001","0000000010100000","1111111111111101","1111111101101001","1111111111010111","0000000001100001","0000000000100110","1111111110100000","1111111101011000","1111111101000100","1111111110100011","0000000001110001","0000000001111011","1111111101001011","1111111010010000","1111111100110100","1111111111100011","0000000001001010","0000000110001110","0000001010011001","0000000110000110","0000000000101101","0000000011000100","0000000100000010","1111111100111111","1111111010101001","0000000001111000","0000000011100000","1111111011110011","1111111001101010","0000000000001001","0000000101000011","0000000111000111","0000000111111001","0000000011001000","1111111110011100","0000000011010100","0000000111010101","1111111111100100","1111111010100110","0000000010011010","0000000101000100","1111111011101000","1111111001010100","0000000001100001","0000000010110100","1111111110011111","0000000001001010","0000000011100111","1111111110110001","1111111111000001","0000000101101001","0000000011010100","1111111100011111","0000000001011100","0000001001010001","0000000100111001","1111111111100110","0000000100111101","0000001001001010","0000000100010000","1111111111001101","1111111110010101","1111111111011001","0000000100100110","0000001010111000","0000001001101111","0000000100100111","0000000011101010","0000000010010001","1111111011111001","1111111000001011","1111111011000110","1111111111010111","0000000010110110","0000000100111000","0000000001100001","1111111011000010","1111111000011000","1111111001110100","1111111101001111","0000000001111101","0000000001110101","1111111010110001","1111111001001010","0000000010000100","0000000110111010","0000000001000111","1111111101000110","1111111111111110","0000000010000001","0000000001101101","0000000010111101","0000000100100110","0000000011011101","1111111110000010","1111110111111100","1111111011101100","0000001000001111","0000001010000001","1111111110111111","1111111110010110","0000000111011010","0000000000011010","1111110001010011","1111111001001100","0000001101010001","0000001011110101","1111111011000111","1111110110011110","1111111110001101","0000000100011000","0000000101011001","0000000001011010","1111111011111100","1111111101001000","0000000010111101","0000000100001101","0000000001111100","0000000000100101","1111111111000011","1111111111100011","0000000001101110","1111111100001010","1111110010110010","1111110101111110","1111111111100000","1111111101011001","1111111001100001","0000000010111000","0000001010010100","0000000100010100","0000000000110010","0000000011111001","1111111111101110","1111111011000001","0000000011000011","0000001000111010","0000000000110001","1111111100111001","0000000101011101","0000000111111000","1111111111111010","1111111101010000","0000000000101000","1111111111110110","1111111110011010","0000000010010010","0000000101011010","0000000011001010","1111111111101001","1111111110111010","0000000001110101","0000000110000000","0000000101100100","1111111111101111","1111111010110101","1111111001100000","1111111010001000","1111111101001110","1111111111110010","1111111011111110","1111110110101000","1111111001000010","1111111111101011","0000000010111100","0000000100001000","0000000100000001","1111111111110011","1111111100000000","1111111101000111","1111111101101011","1111111011100111","1111111101100100","0000000011010001","0000000101010100","0000000010001110","1111111101011001","1111111011011100","0000000001011001","0000001000001010","0000000000111101","1111110011001101","1111110110001101","0000000110010001","0000001010010010","0000000001111011","0000000000101101","0000000110011011","0000000101011010","0000000000001001","0000000001001011","0000000101011011","0000000100010010","0000000000011000","0000000001000001","0000000011001011","1111111110100001","1111110110100101","1111110110101001","1111111101110001","0000000000100100","1111111100010101","1111111000000101","1111111000101000","1111111101101100","0000000010010010","0000000000001100","1111111010110111","1111111010111101","1111111100110011","1111111001100110","1111111000110011","1111111110010100","1111111101101101","1111110101011011","1111110101000000","1111111100101000","1111111101111010","1111111010101100","1111111101100110","0000000010001110","0000000001011010","0000000000010111","0000000100001011","0000001001001001","0000001001000110","0000000000111011","1111110110011000","1111110100011000","1111111001110100","1111111011111110","1111111011001101","1111111101110101","1111111111111001","1111111110011110","1111111111001111","0000000000001100","1111111100111110","1111111111000001","0000001000110011","0000001000100100","1111111011100100","1111110111011001","1111111111110000","0000000010111001","0000000001000011","0000000110100111","0000001100010011","0000000110110011","1111111110110010","1111111101011100","1111111101010010","1111111011000010","1111111011000011","1111111110010000","0000000010000001","0000000011110100","0000000001111111","0000000001001010","0000000110010110","0000001001000101","0000000001010011","1111111010011011","1111111110110011","0000000100010011","0000000100101111","0000001001000110","0000001111000101","0000001010100100","0000000001110010","0000000001100000","0000000011100110","0000000001100011","0000000011101101","0000001000110000","0000000011010000","1111110111101110","1111110110101111","1111111101111111","0000000000110011","0000000000001101","0000000000110001","1111111110111001","1111111100001110","1111111110101000","1111111111101000","1111111000000001","1111110011111000","1111111101100010","0000000101110001","1111111111000010","1111111001001010","0000000010110100","0000001100100000","0000000110110111","1111111110010011","1111111111110010","0000000011001001","0000000001011000","0000000000000001","1111111111111000","1111111101101011","1111111101110101","0000000001101111","0000000001010100","1111111100001001","1111111010101011","1111111100101001","1111111101111001","0000000001111000","0000000110101001","0000000010000110","1111111001000011","1111111011011111","0000000101101100","0000000110001000","1111111110010110","1111111101100010","0000000010111000","0000000001110101","1111111010101010","1111111000010110","1111111100110101","1111111111111001","1111111110110101","1111111111111100","0000000100011010","0000000100011111","1111111111110110","0000000000101111","0000000110001101","0000000001111100","1111110101110000","1111110100111010","0000000000000011","0000000011101011","1111111101010010","1111111100010000","0000000000110000","1111111110011000","1111110111011110","1111110110111111","1111111011111011","1111111111010111","0000000000100001","0000000000000110","1111111110001100","1111111101111110","0000000001010000","0000000100110001","0000000101001010","0000000010000111","1111111110011011","1111111110010110","0000000000101111","1111111111001100","1111111010011011","1111111001011011","1111111010010100","1111110111110110","1111111000111101","0000000010011000","0000000110011010","1111111101000001","1111110110011110","1111111110011001","0000000110101010","0000000011011001","1111111111011001","0000000100001110","0000001000100001","0000000011010010","1111111011100110","1111111011100011","0000000001010010","0000000100100011","0000000010100011","1111111110111000","1111111100011010","1111111011011011","1111111101001101","0000000010000110","0000000100010101","1111111110110010","1111111000000000","1111111001101011","1111111111010100","1111111110011010","1111111010011011","1111111011101010","1111111100110010","1111110111101000","1111110100110110","1111111010101101","0000000001011111","0000000100110111","0000000111011011","0000000100111011","1111111101000111","1111111101000110","0000000101100111","0000000101111111","1111111111101010","0000000010100101","0000000110011100","1111111011000110","1111101110111010","1111110011001011","1111111010111010","1111111011010101","1111111110111100","0000000100110001","0000000001011100","1111111101011110","0000000010001011","0000000010111000","1111111100011110","1111111111000000","0000001000011000","0000001001000001","0000000110001110","0000001000110000","0000000110011110","1111111110011100","1111111110111001","0000000011010101","1111111110001001","1111111000110010","1111111101010111","1111111110101110","1111110111111100","1111111001011100","0000000100111111","0000001000101101","0000000001011000","1111111101110110","0000000100000000","0000001001110000","0000000101001001","1111111010000110","1111110101101011","1111111011010010","0000000010001100","0000000111001100","0000001100000100","0000001011000000","0000000010011000","1111111110011011","0000000010101110","0000000011110110","0000000001000011","0000000011100000","0000000111000010","0000000011010101","1111111101011000","1111111010101101","1111111010010110","1111111111110100","0000001011001000","0000001111100111","0000000111111010","1111111111101011","1111111101111111","1111111110000110","1111111110101000","0000000010000001","0000000101111101","0000000110001111","0000000001110110","1111111100010111","1111111101011101","0000000110001010","0000001011001011","0000000110100100","0000000000101101","1111111110010000","1111111011100001","1111111011010101","0000000000001100","0000000001011100","1111111101010100","1111111110110011","0000000011111001","0000000000000011","1111111001101110","1111111100111000","1111111110010011","1111110101011101","1111110100001100","0000000000101111","0000000011111111","1111111000010000","1111110101100010","0000000000100100","0000000100110110","1111111111100111","1111111111011000","0000000100010001","0000000110000001","0000000100100011","0000000000001100","1111111001110111","1111111001010100","1111111101101001","1111111011001001","1111110100111100","1111111000110111","0000000010011000","0000000100011100","0000000010101100","0000000100000101","0000000100010101","0000000001111111","0000000000101000","1111111110010111","1111111011101100","1111111101100111","1111111111111010","1111111101101000","1111111110011110","0000000100101011","0000000101001001","1111111111101001","1111111110000000","1111111101110001","1111111011011100","1111111111101000","0000000111111000","0000000101101101","1111111110100001","0000000001000000","0000000011110111","1111111010100011","1111110011100101","1111111100100011","0000000111011010","0000000101100000","1111111101110000","1111111100010010","0000000010110001","0000001001100110","0000000111011100","1111111110111001","1111111101001010","0000000010011001","0000000000101000","1111111000110010","1111111001111100","0000000011000001","0000000110110100","0000000101101110","0000000101011011","0000000001110000","1111111100000100","1111111110111111","0000000111000000","0000000110110001","0000000001111101","0000000010111010","0000000011110100","1111111111001010","1111111110101011","0000000100000011","0000000010000011","1111111000100000","1111110110011010","1111111110110111","0000000111001011","0000001000111100","0000000110000101","0000000100111001","0000001000101010","0000001000011110","1111111101111100","1111111000111000","0000000101001011","0000001110101100","0000000110000101","1111111111010101","0000000110010011","0000000110011110","1111111010010111","1111111000001000","0000000001010110","0000000001110010","1111111010101011","1111111011010001","1111111111011110","1111111101100011","1111111011110011","0000000000011100","0000000100010001","0000000001000001","1111111011000011","1111111010000010","1111111111011101","0000000100011011","0000000010111000","1111111110100111","1111111101101010","1111111111000100","0000000000110011","0000000011110000","0000000101101110","0000000010010011","1111111010011110","1111110101000011","1111111000010101","0000000001001110","0000000011100000","1111111100101010","1111111011010001","0000000011100110","0000000100110101","1111111010010101","1111110101110101","1111111100111101","0000000010101101","0000000011111000","0000000110011100","0000000111000011","0000000001111100","1111111101111011","0000000000011010","0000000101010111","0000000101101110","1111111110111110","1111111010000000","0000000001001001","0000001010010101","0000000101001011","1111111011011010","1111111110100111","0000000101111110","0000000100110001","0000000011010001","0000000101000110","0000000001010000","1111111101110000","0000000100101110","0000001010010110","0000000101000100","0000000000110100","0000000010000001","1111111110101100","1111111001010001","1111111001111101","1111111100011001","1111111110010011","0000000011000111","0000000011100101","1111111100011000","1111111100010011","0000000110000111","0000000111100010","1111111111010001","1111111101111000","0000000001111010","0000000000101001","1111111111110101","0000000011000000","0000000000010101","1111111011010101","0000000001000101","0000001000000010","0000000000011110","1111110110111111","1111111101001000","0000000111000010","0000000011100000","1111111010111111","1111111011101000","0000000000100110","0000000000101110","1111111111001011","0000000000011000","0000000000111100","1111111111001001","1111111110101111","0000000000011110","0000000001100110","0000000001100100","1111111111101101","1111111011000100","1111111000010001","1111111010101001","1111111100000001","1111111010110011","1111111111111111","0000001000111011","0000000111000101","1111111111000110","0000000001100001","0000000111001111","0000000001100011","1111111011100001","0000000000100010","0000000010011101","1111111010100011","1111111000101110","0000000000000001","0000000010101011","0000000000010001","0000000000010101","0000000001000110","0000000010011110","0000000110000010","0000000100101110","0000000000000000","0000000100010010","0000001010101011","0000000100000100","1111111101011101","0000000101010001","0000001001010101","1111111111100101","1111111101010101","0000000110110001","0000000110110001","1111111111010101","0000000001011000","0000000101010010","1111111111110010","1111111010100001","1111111001011111","1111110101010000","1111110011110111","1111111100011000","0000000011110101","0000000100001010","0000000101010110","0000000101101000","1111111111000010","1111111010101010","1111111110000110","1111111110110001","1111111010110111","1111111100111010","0000000011000001","0000000011100110","0000000001000011","0000000000101000","1111111111100101","1111111101111101","1111111111100000","0000000000111001","1111111101111000","1111111100000001","0000000001100000","0000001001010010","0000001000111111","1111111111111010","1111111010001011","0000000000000001","0000000111110100","0000000101011100","1111111110100110","1111111101111111","1111111111101111","1111111101100000","1111111011111101","1111111110010111","0000000000110011","0000000010001000","0000000001100110","1111111100011100","1111111010000010","0000000011010101","0000001101010100","0000001010100001","0000000101001000","0000000110100111","0000000010100010","1111110101110110","1111110010110110","1111111011110010","1111111110111110","1111111010101000","1111111001110101","1111111011101011","1111111101000101","0000000001010110","0000000011000101","1111111101010011","1111111011110001","0000000011010110","0000000101000000","1111111111011100","0000000011011101","0000001101010100","0000001001111011","1111111110010010","1111111101000101","0000000011111111","0000000101111100","0000000010100101","1111111110101101","1111111011011101","1111111011111010","0000000001110001","0000000110011001","0000000011101110","1111111101100101","1111111011001111","1111111100111111","1111111101000000","1111111001110110","1111111001101101","1111111110110001","0000000010001000","0000000000110011","0000000000100010","0000000011000001","0000000100000100","0000000011010000","0000000010100111","0000000001100011","0000000000101101","0000000000111001","0000000000010110","0000000001001101","0000000110000110","0000000111001001","1111111111011111","1111111011110111","0000000010110001","0000000100111110","1111111011101111","1111110110010010","1111111010111010","1111111111000100","1111111111111110","0000000010000101","0000000010010000","1111111110101101","1111111100111100","1111111110000001","1111111111100100","0000000010100100","0000000100011100","0000000000110011","1111111100001000","1111111011001110","1111111011000001","1111111011011001","1111111101101001","1111111011101111","1111110111011110","1111111101010010","0000001000011011","0000000111010001","1111111110010101","1111111101000110","1111111111001000","1111111101001110","1111111110111001","0000000010111110","1111111111000000","1111111000100111","1111111010000101","1111111110001100","0000000000010010","0000000010000111","1111111110011010","1111110110100001","1111111000111000","0000000010100100","0000000010000110","1111111101110110","0000000100110101","0000001010111010","0000000100011010","0000000001001101","0000001000110001","0000001010010010","0000000001000100","1111111010111100","1111111100010000","0000000000011001","0000000101000101","0000000100101011","1111111100101000","1111111000100100","0000000000100000","0000001001011100","0000000111100001","1111111110010001","1111110111111110","1111111001011001","1111111110001000","1111111110011001","1111111011010000","1111111100011001","0000000000101010","0000000001101101","0000000010100111");
signal sdatad : array_data:=
--(others=>(others=>'0'));
("0000000000000000","0000001000001101","0000010000010010","0000011000000110","0000011111100000","0000100110011001","0000101100101001","0000110010001010","0000110110110110","0000111010101000","0000111101011011","0000111111001110","0000111111111110","0000111111101010","0000111110010011","0000111011111010","0000111000100001","0000110100001101","0000101111000001","0000101001000100","0000100010011011","0000011011001110","0000010011100100","0000001011100101","0000000011011010","1111111011001011","1111110011000001","1111101011000110","1111100011100000","1111011100011000","1111010101110110","1111010000000001","1111001010111111","1111000110110100","1111000011100110","1111000001011000","1111000000001101","1111000000000100","1111000001000000","1111000010111110","1111000101111101","1111001001111001","1111001110101110","1111010100011000","1111011010101111","1111100001101110","1111101001001110","1111110001000101","1111111001001100","0000000001011010","0000001001100111","0000010001101001","0000011001011001","0000100000101110","0000100111100001","0000101101101001","0000110011000001","0000110111100100","0000111011001011","0000111101110100","0000111111011011","0000111111111111","0000111111100000","0000111101111101","0000111011011001","0000110111110110","0000110011010111","0000101110000011","0000100111111110","0000100001001110","0000011001111010","0000010010001101","0000001010001100","0000000001111111","1111111001110000","1111110001101001","1111101001110001","1111100010001111","1111011011001100","1111010100110011","1111001111001000","1111001010001101","1111000110001010","1111000011001001","1111000001001001","1111000000000111","1111000000000111","1111000001010000","1111000011011101","1111000110100101","1111001010100110","1111001111101000","1111010101011111","1111011011111011","1111100010111001","1111101010100001","1111110010100011","1111111010101000","0000000010101101","0000001010111110","0000010011001000","0000011010101110","0000100001110010","0000101000100101","0000101110110011","0000110011111011","0000111000000011","0000111011101001","0000111110011001","0000111111101010","0000111111101110","0000111111001111","0000111101111010","0000111010111100","0000110110110001","0000110010011010","0000101101100000","0000100110111110","0000011111011101","0000011000011111","0000010001100011","0000001000111110","1111111111101000","1111111000000111","1111110001110001","1111101000110010","1111011100110010","1111010010110001","1111001101110100","1111001010100010","1111000101010100","1111000000111110","1111000010010100","1111000111100010","1111001001110011","1111000110010011","1111000000111100","1110111110101001","1111000000111010","1111000111001100","1111001111110100","1111010111101011","1111011100111100","1111100010110011","1111101101111001","1111111100011011","0000000110100111","0000001001000100","0000001010000000","0000010000110011","0000011100010100","0000100110000000","0000101011010110","0000101110111000","0000110001101110","0000110010100000","0000110010110001","0000110111000101","0000111111011000","0001000100101101","0001000010010101","0000111100100011","0000111001111110","0000111001011110","0000110100110010","0000101010111010","0000100001001101","0000011010011010","0000010011011000","0000001010011011","0000000011001111","1111111111110010","1111111011010100","1111110001100101","1111100110101011","1111100001010111","1111100000000000","1111011010110111","1111010000110100","1111001001101111","1111001001101101","1111001001100000","1111000001101000","1110110110100111","1110110011010111","1110111001111000","1111000001110110","1111000101100001","1111001000100010","1111001111111011","1111011010001010","1111100010100000","1111100111111101","1111101101001100","1111110100100001","1111111110011001","0000001001011010","0000010010010001","0000010110101001","0000011001010000","0000011111001111","0000101000100101","0000101111101010","0000110010001000","0000110100100000","0000111010010101","0001000000000000","0001000000110111","0000111110100000","0000111101010011","0000111101011101","0000111100001000","0000111000010111","0000110010110110","0000101011011011","0000100010010101","0000011001100011","0000010010001000","0000001010110011","0000000011001000","1111111100011101","1111110110001111","1111101110000010","1111100100110011","1111011110010111","1111011001110110","1111010001110000","1111000110011100","1111000000011000","1111000011001101","1111000110110110","1111000011111001","1110111110111011","1110111111110011","1111000100111000","1111000111110111","1111001001011110","1111001110010100","1111010100110110","1111011000100100","1111011011111001","1111100100100011","1111110000010101","1111110111110100","1111111011011001","0000000010101011","0000001111000110","0000011001001101","0000011101010000","0000100000111111","0000101001101000","0000110100000010","0000111010110110","0000111101111100","0000111111111011","0001000001010010","0001000001001111","0000111111110101","0000111100101001","0000110111001110","0000110010000000","0000110000010111","0000110000110101","0000101101111101","0000100110001011","0000011101110011","0000010111011110","0000010000001011","0000000101001110","1111111001000111","1111101111101011","1111101001010010","1111100100100010","1111100000100110","1111011011110111","1111010100100011","1111001100010110","1111000111100000","1111000110011010","1111000100100110","1110111111101100","1110111011010110","1110111011111010","1111000001011111","1111001001101000","1111010001111010","1111010111101000","1111011001011110","1111011010100111","1111011111011111","1111100111010010","1111101101101000","1111110010100111","1111111010101001","0000000101110010","0000001110111011","0000010101001011","0000011101101000","0000101001011111","0000110010010001","0000110011110001","0000110010100001","0000110100000001","0000110111011110","0000111010001010","0000111100011000","0000111110001001","0000111101000100","0000111001100100","0000110111111101","0000111000010111","0000110100011000","0000101001001111","0000011101111010","0000011001001010","0000010111110010","0000010010010001","0000000111101000","1111111100011010","1111110011001011","1111101011010000","1111100100001000","1111011101010010","1111010101011110","1111001101100000","1111001000110111","1111001000010000","1111000111110101","1111000101000111","1111000010001101","1111000001000000","1111000000010110","1111000000111011","1111000101111101","1111001101110101","1111010001011010","1111001111101010","1111010001110110","1111011101111001","1111101100001001","1111110011001001","1111110110001100","1111111110001000","0000001001101110","0000010001001100","0000010101000111","0000011101010000","0000101001110100","0000110010100011","0000110101000000","0000110111101100","0000111101111010","0001000011000011","0001000100101010","0001000110101110","0001001010001100","0001001001000111","0001000000110010","0000110111001111","0000110001110110","0000101110000110","0000101000001100","0000100001101101","0000011100110011","0000010111010001","0000001111001000","0000000110110001","1111111111110011","1111110111101011","1111101101000011","1111100011011001","1111011101000010","1111010111000110","1111001111000000","1111000111011100","1111000011110111","1111000011011000","1111000011011001","1111000011001101","1111000010011110","1111000000100011","1110111111100010","1111000010111001","1111001001100111","1111001111000010","1111010011000010","1111011010011011","1111100101101011","1111101110110011","1111110011011101","1111111001001110","0000000011110110","0000001110100110","0000010100100110","0000011000100011","0000011111000110","0000100111001111","0000101101101100","0000110010101010","0000110110110011","0000110111111001","0000110101111111","0000110110110111","0000111110010111","0001000111000110","0001001000100011","0001000001010101","0000110110101111","0000101101010110","0000100110101000","0000100010101111","0000011111101100","0000011001011101","0000001110111111","0000000100100000","1111111101010000","1111110111000000","1111101111011000","1111101001001011","1111100110011100","1111100010010011","1111010111101101","1111001011000001","1111000100101111","1111000100101011","1111000010111011","1110111101011011","1110111011001111","1111000000011101","1111000111001000","1111001000011011","1111000110100011","1111001000101100","1111010001000000","1111011011011010","1111100011101110","1111101001001011","1111101101100111","1111110011101110","1111111100110001","0000000110110011","0000001110111100","0000010101101001","0000011101100000","0000100101101101","0000101010011100","0000101100001000","0000110000010011","0000111000100100","0000111110111111","0000111111000100","0000111100111010","0000111110001011","0001000000111000","0000111111101111","0000111011000001","0000110110110111","0000110011010011","0000101101011110","0000100110010110","0000100001011001","0000011101101111","0000010111001001","0000001101001001","0000000010101000","1111110111101000","1111101010011001","1111011101111000","1111010111011100","1111010101110010","1111010001110110","1111001010000110","1111000100110011","1111000100100110","1111000011011111","1110111101100111","1110111001010100","1110111101101100","1111000110110001","1111001010111011","1111001000101001","1111000111000011","1111001010111100","1111010010110010","1111011100110001","1111101000111101","1111110100010100","1111111001101110","1111111010110100","0000000000101000","0000001110101011","0000011011111100","0000011111000111","0000011100111011","0000100001101100","0000101111000010","0000111001110010","0000111010101001","0000111000000111","0000111011100110","0001000011110111","0001001000000111","0001000100101011","0000111110001010","0000111001100111","0000110110110111","0000110010101001","0000101010101110","0000011111100110","0000010100110001","0000001110011000","0000001100010000","0000001000110011","0000000000001010","1111110110010100","1111110001011111","1111101111100000","1111100111110010","1111011000111100","1111001100101111","1111001010100100","1111001100100100","1111001001001110","1111000010000101","1111000000010101","1111000101001110","1111001000000000","1111000100001101","1111000000100111","1111000100011110","1111001101100100","1111010101110111","1111011100100011","1111100011111000","1111101010101010","1111101110101001","1111110010001100","1111111001101011","0000000100100011","0000001110000101","0000010100011110","0000011010110000","0000100011100101","0000101101001001","0000110011010000","0000110100011001","0000110011111011","0000110110101100","0000111100111000","0001000001010011","0001000000001011","0000111100000001","0000111000011000","0000110011111001","0000101101010100","0000101001010111","0000101011000101","0000101010010110","0000011101110111","0000001100001110","0000000100110110","0000000111111000","0000000101000101","1111110101101100","1111100110011001","1111100001000010","1111011101101111","1111010100010111","1111001100000001","1111001100001111","1111001100111101","1111000100111000","1110111011101110","1110111101011111","1111000101000011","1111000101000100","1110111110111101","1110111111000101","1111000110111101","1111001101010100","1111010000110000","1111011000101010","1111100100100100","1111101011100001","1111101100101010","1111110001010011","1111111100101110","0000000111101101","0000001110001100","0000010100100111","0000011101111000","0000100111011100","0000110000100000","0000111001111000","0000111110110101","0000111010011001","0000110011011010","0000110101110000","0000111110110111","0001000000010000","0000110111000111","0000110001000111","0000110101100010","0000111001110001","0000110011110001","0000101001000101","0000100010001110","0000011100000011","0000010000100010","0000000011110011","1111111101000000","1111111001111100","1111110011110101","1111101010111111","1111100100000100","1111011111000001","1111011000101110","1111010001100111","1111001011101000","1111000101011101","1110111110001110","1110111001101111","1110111010111100","1110111110101100","1111000000111111","1111000011000100","1111000111001011","1111001011101100","1111001111111000","1111010111110001","1111100100110000","1111101111111001","1111110010110011","1111110010000101","1111110111000010","0000000010010110","0000001100110010","0000010010111001","0000011000100011","0000100001001111","0000101011000101","0000110010001001","0000110100011110","0000110011010001","0000110010101110","0000110111000110","0000111111000101","0001000011110011","0001000001000110","0000111010110010","0000110110011101","0000110100001001","0000110001011000","0000101110111011","0000101101111000","0000101010100110","0000100001000011","0000010100000110","0000001001111100","0000000010111111","1111111010100001","1111101111010111","1111100101011110","1111011111001001","1111011010010011","1111010100111101","1111001111100101","1111001010100111","1111000110000100","1111000011001000","1111000010000011","1110111111011101","1110111000110111","1110110011001100","1110110110101001","1111000011001010","1111001111011011","1111010100110000","1111010110100000","1111011011010101","1111100100011010","1111101110010100","1111110110011111","1111111100100001","0000000000111101","0000000110000010","0000001110101110","0000011010100111","0000100100110010","0000101001100111","0000101011110100","0000110000101101","0000111000101111","0000111110111111","0001000000000000","0000111110010011","0000111110010001","0000111111111000","0000111110111001","0000111001010011","0000110010001111","0000101100111110","0000100111110001","0000100000000001","0000011001000111","0000011000101110","0000011011111101","0000010111010100","0000000101011111","1111110000001100","1111100100110011","1111100100000111","1111100011100001","1111011011111010","1111010000110011","1111001001000011","1111000110100010","1111000110001011","1111000100011110","1111000000100011","1110111100110011","1110111100110111","1111000001010111","1111000110100100","1111001001000100","1111001010011101","1111001110110001","1111010110011100","1111011101111101","1111100011000011","1111100111100111","1111101110111101","1111111001110111","0000000101101101","0000001110111110","0000010101000001","0000011010111100","0000100011100000","0000101100111000","0000110010101111","0000110100100000","0000110101111111","0000111001011000","0000111100100110","0000111110011111","0001000001110100","0001000111011000","0001001001001110","0001000001001010","0000110010101000","0000101000000001","0000100101110001","0000100101011011","0000011111100011","0000010101011101","0000001101001010","0000000110111111","1111111101111011","1111110001100000","1111101000010001","1111100101110010","1111100100100001","1111011110010101","1111010110000101","1111010010001111","1111010001101010","1111001101100000","1111000101010100","1111000000010010","1111000001110101","1111000100110001","1111000100011101","1111000011110000","1111000111000011","1111001101010000","1111010010110110","1111010111000111","1111011010111010","1111011110010000","1111100010101000","1111101011101011","1111111001111100","0000001000100000","0000010010100100","0000011000000000","0000011010110010","0000011100100100","0000100000110101","0000101011011111","0000111001111110","0001000011010001","0001000011000101","0000111111100000","0000111111011010","0001000000110000","0000111110010111","0000111001101011","0000110111011000","0000110110001010","0000110000100100","0000100110110101","0000011110111011","0000011011011000","0000011000010000","0000010001111110","0000001001010111","1111111111111010","1111110101110111","1111101101000000","1111100111111110","1111100101000111","1111011110111110","1111010100010101","1111001010111101","1111000111001100","1111000101101111","1111000001110101","1110111101011100","1110111101101101","1111000001110100","1111000011111111","1111000010101111","1111000010111001","1111001000000011","1111010000011000","1111011001000101","1111100010000100","1111101011001101","1111110010010101","1111110110110110","1111111011100100","0000000010101010","0000001010111000","0000010010110101","0000011011110010","0000100110001010","0000101110110010","0000110010111101","0000110101000000","0000111000101100","0000111101100000","0001000000001100","0001000000100011","0001000001000111","0001000001101100","0000111110100100","0000110110011100","0000101110000001","0000101011000001","0000101100101010","0000101011010110","0000100000110100","0000010000000110","0000000011001011","1111111111010000","1111111101111110","1111110101110000","1111100111011100","1111011101011011","1111011100001100","1111011011000101","1111010001001011","1111000011100000","1110111110001000","1111000010100000","1111000101111011","1111000010000011","1110111101011110","1111000000000100","1111000110111101","1111001001110111","1111000111110100","1111000111011100","1111001101010011","1111010111011100","1111100001110101","1111101010011110","1111110001011011","1111111000011010","0000000001101000","0000001100010000","0000010100000111","0000011000010010","0000011110011010","0000101010011000","0000110110001011","0000111001011111","0000110110110000","0000111000000011","0000111111100000","0001000100101001","0001000010000100","0000111100101111","0000111010011110","0000111001110101","0000110111101001","0000110101000001","0000110010110001","0000101101010011","0000100010100010","0000010110100101","0000001101100011","0000000101101011","1111111100010110","1111110011110110","1111101110111111","1111101011100000","1111100101111110","1111011111011110","1111011010101000","1111010110011101","1111010000100100","1111001001101100","1111000011110100","1110111110110001","1110111010100100","1110111001111101","1110111110101010","1111000101011101","1111001001110110","1111001011111011","1111001111001101","1111010101001111","1111011100001110","1111100010011000","1111101000010000","1111101111110001","1111111001111000","0000000100101100","0000001101001000","0000010011010010","0000011011000010","0000100101111110","0000101111100000","0000110011000100","0000110011100000","0000110110110001","0000111100011010","0000111111000000","0000111101110110","0000111101100110","0000111110111111","0000111100111001","0000110101110010","0000101111110011","0000101111010111","0000101111111000","0000101010011011","0000011111100010","0000010101011100","0000001110111010","0000001001001010","0000000001011100","1111111000110001","1111110000111010","1111101001000110","1111011111111001","1111010110111110","1111010001110111","1111010000100011","1111001110000111","1111000111001110","1110111111101000","1110111101010111","1111000000010010","1111000010111111","1111000011001100","1111000011110010","1111000110111011","1111001011110111","1111010010011110","1111011010111101","1111100001111111","1111100100100101","1111100111010001","1111110001010100");
--("1111111111111111","0000001000001101","0000010000010010","0000011000000110","0000011111100000","0000100110011001","0000101100101001","0000110010001010","0000110110110110","0000111010101000","0000111101011011","0000111111001110","0000111111111110","0000111111101010","0000111110010011","0000111011111010","0000111000100001","0000110100001101","0000101111000001","0000101001000100","0000100010011011","0000011011001110","0000010011100100","0000001011100101","0000000011011010","1111111011001011","1111110011000001","1111101011000110","1111100011100000","1111011100011000","1111010101110110","1111010000000001","1111001010111111","1111000110110100","1111000011100110","1111000001011000","1111000000001101","1111000000000100","1111000001000000","1111000010111110","1111000101111101","1111001001111001","1111001110101110","1111010100011000","1111011010101111","1111100001101110","1111101001001110","1111110001000101","1111111001001100","0000000001011010","0000001001100111","0000010001101001","0000011001011001","0000100000101110","0000100111100001","0000101101101001","0000110011000001","0000110111100100","0000111011001011","0000111101110100","0000111111011011","0000111111111111","0000111111100000","0000111101111101","0000111011011001","0000110111110110","0000110011010111","0000101110000011","0000100111111110","0000100001001110","0000011001111011","0000010010001101","0000001010001100","0000000001111111","1111111001110000","1111110001101001","1111101001110001","1111100010001111","1111011011001101","1111010100110011","1111001111000111","1111001010001101","1111000110001011","1111000011001001","1111000001001000","1111000000000111","1111000000000111","1111000001010000","1111000011011101","1111000110100101","1111001010100111","1111001111101000","1111010101011110","1111011011111011","1111100010111010","1111101010100001","1111110010100010","1111111010100111","0000000010101111","0000001010111110","0000010011000111","0000011010101110","0000100001110011","0000101000100101","0000101110110001","0000110011111010","0000111000000101","0000111011101001","0000111110010111","0000111111101010","0000111111110000","0000111111010000","0000111101110110","0000111010111011","0000110110110101","0000110010011100","0000101101011010","0000100110111100","0000011111100110","0000011000100010","0000010001010110","0000001000111001","1111111111111110","1111111000010000","1111110001000011","1111101000011101","1111100000000001","1111011011100110","1111011010110011","1111010111101101","1111001110110111","1111000100100011","1110111111010101","1111000000000111","1111000010100000","1111000010110111","1111000001000010","1110111110111001","1110111111011000","1111000100111011","1111001110100000","1111010111010110","1111011100001101","1111011111100111","1111100110001111","1111110000110010","1111111100011001","0000000111011110","0000010010100110","0000011101001100","0000100100110101","0000101000100110","0000101010110010","0000101110001001","0000110011100000","0000111010000001","0000111111111001","0001000010110110","0001000010001010","0001000000100000","0001000000111110","0001000010000010","0000111111000010","0000110111100010","0000110001000011","0000101110010110","0000101010010011","0000011111110110","0000010011001110","0000001100001101","0000001001110001","0000000011101101","1111111000000101","1111101110010011","1111101010100110","1111100111110010","1111100001001100","1111011010001001","1111010110001100","1111010001010111","1111000111110011","1110111110011101","1110111100001111","1110111110111101","1110111111111101","1110111111100011","1111000010111011","1111001001110100","1111001111000110","1111010010001101","1111010111001001","1111011110011100","1111100101001101","1111101100000000","1111110101100001","1111111111011011","0000000101011011","0000001010010101","0000010100100101","0000100010001011","0000101010001101","0000101011011000","0000101110001101","0000110110101010","0000111110001010","0000111111100001","0000111110111011","0001000000111010","0001000010011001","0000111111100000","0000111011000001","0000111000110101","0000110111000000","0000110001111010","0000101010001101","0000100010011100","0000011011000111","0000010100111001","0000010001001000","0000001101000010","0000000011010101","1111110101100101","1111101100011111","1111101010010101","1111100101111100","1111011001000101","1111001011011100","1111000110110011","1111000111110110","1111000100111000","1110111110000000","1110111011100101","1110111111101011","1111000011111110","1111000101010011","1111000110111011","1111001010011101","1111001101101011","1111010001001001","1111011000011101","1111100010001101","1111101000100100","1111101011101000","1111110010101000","1111111111101110","0000001011000010","0000001111001011","0000010010100100","0000011101011000","0000101100010000","0000110101100101","0000110111101011","0000111000101010","0000111010110100","0000111011000011","0000111010000001","0000111100101111","0001000010010011","0001000010111101","0000111100101010","0000110111010110","0000110111011111","0000110101110010","0000101011100100","0000011111000000","0000011001010111","0000010111001111","0000001110010001","1111111110111000","1111110100001110","1111110010111001","1111110010110011","1111101100011000","1111100001110111","1111011001000011","1111010011010000","1111001111000101","1111001011110110","1111001000100001","1111000100001011","1111000000111101","1111000010001101","1111000110111101","1111001010110000","1111001011110111","1111001100000101","1111001100100011","1111001101111110","1111010011100101","1111011111001011","1111101011111001","1111110100000000","1111111001111000","0000000011111011","0000010000111000","0000011001100010","0000011101000111","0000100001111000","0000101001001101","0000101101010010","0000101100100011","0000101101100010","0000110011111001","0000111010100011","0000111100110010","0000111101010101","0000111111011001","0000111111111110","0000111011011011","0000110100011100","0000110000001110","0000101111000100","0000101101010111","0000101000101110","0000100000110000","0000010101010110","0000000111100011","1111111010110100","1111110010100011","1111101110101110","1111101011110110","1111100110000100","1111011100111101","1111010100111111","1111010011000101","1111010101011010","1111010011101000","1111001001011010","1110111101011000","1110111001000101","1110111100111101","1111000001110111","1111000011111111","1111000110001001","1111001010111001","1111010001001010","1111010111111011","1111011111100010","1111100110100101","1111101010110101","1111101110000110","1111110101000000","1111111111101011","0000001000111010","0000001110011001","0000010100100101","0000011111001110","0000101010101110","0000110000110000","0000110000111110","0000110001010010","0000110110010011","0000111110000110","0001000010101101","0001000000100101","0000111010100011","0000110111001000","0000111000111010","0000111010111011","0000110110001001","0000101010011010","0000011110111101","0000011001110010","0000011001001101","0000010110111110","0000001111100100","0000000100101000","1111111001100111","1111110000010010","1111101000010111","1111100001001100","1111011010110100","1111010101001101","1111001111011110","1111001000111100","1111000010110011","1110111110111001","1110111100111110","1110111011011101","1110111011011100","1111000000001000","1111001000101001","1111001110111000","1111001111011100","1111001111000111","1111010011100010","1111011010101100","1111011111110100","1111100101001100","1111110000100010","1111111110110011","0000000110000110","0000000101011101","0000001000011001","0000010110001100","0000100110101000","0000101101111111","0000101101011000","0000101110010110","0000110011110100","0000111000011011","0000111001010110","0000111001100001","0000111010011110","0000111001101000","0000110101110110","0000110001110001","0000101111000101","0000101100011100","0000101000110010","0000100100101101","0000011111111101","0000011001100011","0000010010100010","0000001100101011","0000000110100010","1111111101000111","1111110001011111","1111101000100010","1111100100000000","1111011111111100","1111011000011010","1111001110010010","1111000101011011","1111000000011100","1110111111000101","1110111110110001","1110111100111110","1110111010111011","1110111101010011","1111000101101110","1111001110110100","1111010010101001","1111010011001101","1111010111100000","1111100001010110","1111101011011001","1111110001110001","1111110110111111","1111111110110000","0000001000001100","0000010000000101","0000010101110111","0000011011111111","0000100011110000","0000101011000110","0000101111001110","0000110001100101","0000110111110000","0001000011100111","0001001101100000","0001001011111010","0001000001001101","0000111010010011","0000111100110111","0000111110111111","0000110110010010","0000100111111011","0000100000101111","0000100010010001","0000100010010010","0000011010011111","0000001110110100","0000000100001101","1111111011010001","1111110100101000","1111110001011101","1111101101100110","1111100010110000","1111010100010000","1111001110000000","1111010011000101","1111010110111011","1111001110111100","1111000010000000","1110111101001111","1111000000100011","1111000001111000","1110111111101000","1111000010000010","1111001010110001","1111010000110010","1111010000000011","1111010001001110","1111011011100011","1111101001100010","1111110010111001","1111111001001001","0000000001100000","0000001001110101","0000001101101111","0000010001001001","0000011010011110","0000100110011100","0000101100101010","0000101110001110","0000110100000001","0000111110101010","0001000100001011","0000111111110011","0000111001010101","0000111001001010","0000111101100000","0000111111100110","0000111100010100","0000110100100100","0000101010111010","0000100011101010","0000100001011001","0000011111111000","0000011000100000","0000001100110011","0000000100100101","0000000000101011","1111111000101001","1111101001000100","1111011010100001","1111010101011100","1111010110100101","1111010101011011","1111001111100101","1111000111111100","1111000000100010","1110111011100001","1110111100110101","1111000100010010","1111001010010000","1111001000101010","1111000011101110","1111000100000010","1111001010101010","1111010001100110","1111010101101010","1111011001110101","1111100001100010","1111101100011111","1111111000011011","0000000011001010","0000001010111101","0000010000010100","0000010110101111","0000100000101011","0000101011010010","0000110001001011","0000110001100000","0000110001001001","0000110100101001","0000111011001000","0001000000010010","0001000001011000","0000111111001111","0000111100011001","0000111010010010","0000111000011000","0000110101010001","0000110000101100","0000101100000010","0000100111110111","0000100001110100","0000010110110110","0000001000011000","1111111100011100","1111110110110111","1111110100001001","1111101110010010","1111100100111100","1111011100001101","1111010100100100","1111001010100000","1110111111100110","1110111011111101","1111000010001000","1111001000001100","1111000100010100","1110111010111110","1110111000011001","1110111111000111","1111000110110000","1111001010101101","1111001111100100","1111011000000110","1111011111001100","1111100001000001","1111100010011111","1111101001100100","1111110100011110","1111111110010010","0000000111100100","0000010011100110","0000100000000110","0000100111000101","0000101000101011","0000101011111100","0000110100011011","0000111100100010","0000111110100010","0000111110000100","0001000010100010","0001001010000000","0001001010000001","0000111111100110","0000110101111001","0000110110100100","0000111010100010","0000110100001110","0000100100110101","0000011010110000","0000011010101111","0000011000101101","0000001011110111","1111111100111010","1111110111010000","1111110110100010","1111101110111000","1111100000110100","1111010111010111","1111010101010100","1111010001111011","1111001000111010","1111000001010000","1111000000011010","1111000001010011","1110111110010010","1110111011111011","1111000001011101","1111001011100111","1111010000001101","1111001101011000","1111001100111100","1111010110001010","1111100011101010","1111101011011010","1111101100011011","1111101110010101","1111110101111011","0000000000000101","0000001000101000","0000010000000101","0000011000010111","0000100000010100","0000100110000001","0000101010100011","0000110000010101","0000110111010010","0000111101001101","0001000000011011","0001000000100001","0000111110001011","0000111011100000","0000111010010110","0000111000110111","0000110011100001","0000101011110101","0000101000000110","0000101001010100","0000100111011011","0000011100101011","0000001111010111","0000001000100011","0000000101100011","1111111100100001","1111101101101001","1111100100000001","1111100011111010","1111100011101001","1111011011001000","1111010000001000","1111001011001101","1111001001000101","1111000001011011","1110110110101101","1110110011100011","1110111010001111","1111000001111110","1111000100110010","1111000110011100","1111001011101001","1111010011001011","1111011010010001","1111100000011110","1111100101011101","1111101001100111","1111110001101011","0000000001011000","0000010001111010","0000010111100110","0000010011101010","0000010100100011","0000100000010010","0000101011010111","0000101100010001","0000101011001100","0000110011010001","0000111111000101","0001000010001000","0000111101100001","0000111100010100","0000111111111110","0000111111101100","0000111001011000","0000110100100110","0000110100000100","0000110001011111","0000101001111001","0000100010010010","0000011100111110","0000010100101011","0000000110110101","1111111001110100","1111110011100110","1111110000110111","1111101010111111","1111100010000001","1111011010111101","1111010111001001","1111010010010110","1111001001100101","1111000000010000","1110111100101110","1111000000001000","1111000100001101","1111000011001100","1111000000000101","1111000010011010","1111001010110111","1111010010000101","1111010011111100","1111010100110011","1111011001011100","1111100000100001","1111100111111001","1111110001010000","1111111100111000","0000000110000000","0000001010011000","0000001111011001","0000011001101101","0000100101001001","0000101011110011","0000101111011100","0000110100111010","0000111010110111","0000111101011110","0000111110110111","0001000011011010","0001001000100000","0001000111100011","0001000000101100","0000111010010110","0000110111010010","0000110100100101","0000110000010001","0000101010111111","0000100100001010","0000011010110111","0000010001110101","0000001011111011","0000000110000110","1111111011011101","1111101101111110","1111100011100101","1111011100110100","1111010101110110","1111001111010011","1111001100110101","1111001011011100","1111000100000000","1110111000101110","1110110101001110","1110111101001011","1111000101011010","1111000100010011","1110111111111100","1111000011110011","1111001111001111","1111011000100000","1111011100110101","1111100010111101","1111101110000111","1111111000001101","1111111011101111","1111111100001000","0000000000000000","0000001000000101","0000010000100001","0000011000001001","0000100000100011","0000101000111001","0000101110011000","0000110001111111","0000110111111101","0000111111010100","0001000000100011","0000111001000010","0000110010011011","0000110110110011","0001000001010111","0001000100001010","0000111011110111","0000110010101101","0000101110100111","0000101000011101","0000011011001001","0000001111010011","0000001110000110","0000010000011101","0000001000000011","1111110100111000","1111100100111001","1111011111010101","1111011100101110","1111010101100110","1111001101100011","1111001010110101","1111001011100000","1111001001101100","1111000100110110","1111000001000011","1111000000000101","1111000000101100","1111000010100000","1111000110010110","1111001011110110","1111010001110011","1111010111110001","1111011100111101","1111011111101011","1111100000111001","1111100101110110","1111110010001101","0000000001101100","0000001100010001","0000010000100000","0000010100111101","0000011110001001","0000101000010001","0000101101110001","0000101111110001","0000110011011101","0000111001101101","0000111110100101","0000111111111001","0000111111101101","0001000000001011","0001000000101101","0000111111011111","0000111011011110","0000110100111011","0000101110010100","0000101011000010","0000101010001101","0000100101001101","0000010111110110","0000000111100110","1111111101000111","1111111000100011","1111110011000111","1111101010110101","1111100100001101","1111100000011001","1111011010110101","1111010010011111","1111001100101000","1111001010111011","1111000111100111","1111000000001111","1110111011110001","1110111111110001","1111000110100110","1111000111110100","1111000100111000","1111000101100101","1111001100001011","1111010100011101","1111011100010001","1111100101000101","1111101110100010","1111110110000101","1111111011110011","0000000010010111","0000001010110000","0000010011111111","0000011101110010","0000100111010010","0000101100110011","0000101100100101","0000101100000100","0000110010011010","0000111101101101","0001000100001011","0001000001000110","0000111010100111","0000111000011100","0000111010100010","0000111011111101","0000111010001100","0000110101111100","0000101111101010","0000100111101100","0000100000000000","0000011010011001","0000010101101100","0000001111100000","0000000111100100","1111111111001111","1111110111000000","1111101110100000","1111100110001111","1111011111000100","1111011000111010","1111010011100000","1111001111000001","1111001010101001","1111000100101101","1110111110010110","1110111100001000","1111000000000111","1111000101100110","1111000110101100","1111000100100111","1111000101110100","1111001100110110","1111010101100011","1111011011100111","1111011111101100","1111100101000011","1111101101011001","1111110111111000","0000000010000100","0000001001011101","0000001110001100","0000010100000100","0000011110001110","0000101010001100","0000110010100111","0000110110001111","0000111000011111","0000111011010000","0000111100111001","0000111101000110","0000111110101001","0001000001111001","0001000010000111","0000111100000011","0000110011100010","0000101110011101","0000101100010110","0000101000000011","0000011111111010","0000010111010100","0000010000000111","0000000111110001","1111111100111100","1111110011100000","1111110000000011","1111110000111011","1111101111001001","1111100101111111","1111011000001010","1111001100101110","1111000111011110","1111000101011101","1111000001101011","1110111100011100","1110111010111101","1110111110111101","1111000011000110","1111000011000011","1111000010111101","1111001000111100","1111010010001010","1111010110010001","1111010101010100","1111011000111101","1111100110000100","1111110101100010","1111111111001001","0000000100010000","0000001010101010","0000010011100000","0000011100101010","0000100101110101","0000101110001101","0000110010000001","0000110000100001","0000110000000110","0000110101110110","0000111100111111","0000111101111101","0000111010001110","0000111001001000","0000111011100010","0000111011010100","0000110110001110","0000110000101000","0000101100110010","0000100111100110","0000011111100110","0000010111110111","0000010001000110","0000000111000110","1111111001000100","1111101101111001","1111101010100110","1111101001011010","1111100001010000","1111010011101101","1111001011100110","1111001101100001","1111010000111101","1111001100100110","1111000011010100","1110111111000101","1111000010011100","1111000110001111","1111000101100000","1111000011111101","1111000110011011","1111001011011100","1111010000000011","1111010110001110","1111100000100010","1111101011011011","1111110001101100","1111110101010111","1111111100100010","0000000111000011","0000001110110111","0000010010011010","0000010110111011","0000011111011001","0000101000100110","0000101111110011","0000110110001100","0000111011110101","0000111110011111","0000111111010101","0001000010010001","0001000101100100","0001000010111010","0000111011010011","0000111000000010","0000111011010110","0000111010111101","0000110000100011","0000100100101101","0000100000101010","0000011110111011","0000010101011111","0000000110101001","1111111011010110","1111110011110000","1111101010111011","1111100011100100","1111100010011100","1111100001001010","1111010110001011","1111000110111100","1111000001110000","1111000110100011","1111000111001010","1110111111001001","1110111001110100","1110111101100110","1111000010010011","1111000010000000","1111000011010010","1111001011010010","1111010011110100","1111010111110111","1111011101010110","1111101001001110","1111110101010001","1111111011000000","1111111110110100","0000000110101110","0000001111010011","0000010011111111","0000011001000000","0000100011001010","0000101101011010","0000110001001110","0000110010010111","0000110111100011","0000111101011101","0000111100110110","0000111000110111","0000111010111001","0001000010011110","0001000101011001","0000111111011010","0000110110111111","0000110001100011","0000101100100000","0000100100110110","0000011101000100","0000010111111010","0000010010111101","0000001010011110","1111111110110011","1111110011000100","1111101001001110","1111100001011101","1111011011010100","1111010110000001","1111010000111111","1111001100011111","1111001000100000","1111000011110111","1110111110101011","1110111100011111","1111000000000000","1111000101010011","1111000101101100","1111000001111011","1111000011001101","1111001110101010","1111011101010110","1111100101011100","1111100111011011","1111101011011111","1111110100101000","1111111101101110","0000000011100001","0000001001010110","0000010001111100","0000011010100000","0000100000101111","0000100111100000","0000110000101111","0000111000011010","0000111010111110","0000111100000111","0001000000010101","0001000100001000","0001000001010000","0000111010001101","0000110111011101","0000111010010010","0000111010101100","0000110011110111","0000101010100110","0000100100100110","0000100000001111","0000011001000110","0000001111110110","0000001000011101","0000000011011110","1111111101101110","1111110101011110","1111101100010011","1111100011110011","1111011011010000","1111010001111101","1111001010001000","1111000111010001","1111001000111110","1111001001110010","1111000101100011","1110111111100011","1110111110101010","1111000011011101","1111000110111100","1111000100100100","1111000001001010","1111000100100011","1111001111100010","1111011011110001","1111100011111001","1111101000011010","1111101101100010","1111110110010100","0000000001101101","0000001011101110","0000010010001101","0000010111100011","0000011110110100","0000100110110010","0000101100100000","0000110000110100","0000110110010101","0000111011001110","0000111011011100","0000111000111010","0000111010001011","0001000000001000","0001000100011001","0001000010111000","0000111101000000","0000110011010000","0000100101010101","0000011010000011","0000011010111111","0000100011100101","0000100001100011","0000001101101101","1111111000011001","1111110010110110","1111110110111100","1111110010100001","1111100010111110","1111010110000111","1111010011000110","1111010010000100","1111001011101010","1111000011100110","1110111111101110","1110111110101010","1110111100110010","1110111011100000","1110111110100000","1111000101001111","1111001011101011","1111001111100010","1111010010001000","1111010101111001","1111011011110011","1111100011000010","1111101010100011","1111110001111110","1111111000101100","1111111101110010","0000000010101000","0000001011100101","0000011010001010","0000100111111101","0000101101000011","0000101011010000","0000101100001101","0000110011011110","0000111001111111","0000111010001110","0000111001001011","0000111101011010","0001000011110011","0001000100011101","0000111110110111","0000111001011101","0000110110110111","0000110010111010","0000101010000111","0000011110100010","0000010100000100","0000001100010101","0000000111001010","0000000011011100","1111111110001001","1111110100001111","1111100110111111","1111011100000010","1111010111000110","1111010101011000","1111010001100001","1111001011001010","1111000110111110","1111000110111100","1111000110100011","1111000001011110","1110111011101110","1110111101100110","1111000111111100","1111010001110010","1111010011110101","1111010001100010","1111010011010100","1111011011011100","1111100101011010","1111101101100010","1111110100001110","1111111010100111","0000000001000111","0000001000110110","0000010010101110","0000011101000100","0000100101000100","0000101010110111","0000110001000101","0000111000011010","0000111110101011","0001000010001001","0001000011011110","0001000100010101","0001000101011011","0001000101101110","0001000010110100","0000111011011111","0000110010101011","0000101100111110","0000101010011111","0000100110100110","0000011111010110","0000011000000100","0000010010100011","0000001011000111","1111111111110001","1111110101010100","1111101111100101","1111101010010000","1111011111110100","1111010011001110","1111001011000011","1111000111010010","1111000011100001","1110111111101100","1110111110011100","1110111110011110","1110111101110100","1111000000000001","1111000111110010","1111001110011010","1111001100001101","1111000110011101","1111001001010011","1111010101001111","1111011111010101","1111100011101000","1111101010000101","1111110111000110","0000000011101001","0000001001100101","0000001100111010","0000010011011110","0000011011111011","0000100010101011","0000101000110011","0000110000111111","0000111010000001","0001000000011101","0001000010101110","0001000001011110","0000111110101101","0000111101011011","0000111110010000","0000111101100110","0000111000110100","0000110011010101","0000110001100101","0000110001000100","0000101011110111","0000100001110001","0000010111001010","0000001101000100","0000000001101100","1111110111011100","1111110010011011","1111101111111010","1111101000100000","1111011011111100","1111010010010111","1111010000001001","1111010000000000","1111001011011100","1111000011010101","1110111101001000","1110111011101011","1110111101011100","1110111111001001","1110111111000001","1110111110111001","1111000010110010","1111001011101111","1111010101101110","1111011100110101","1111100010001011","1111101000111111","1111110001010000","1111111000110101","1111111111101001","0000000111001100","0000001111001111","0000010110011000","0000011100111011","0000100100010101","0000101100011111","0000110011100110","0000110111111111","0000111001100100","0000111001111101","0000111011010101","0000111101100000","0000111101111101","0000111100101101","0000111101110011","0001000001100011","0000111111110111","0000110010100100","0000100001100100","0000011010100111","0000011101110011","0000011101000010","0000010000011010","0000000000001010","1111110110111110","1111110100000010","1111110000011111","1111101010000011","1111100001111101","1111011000010000","1111001110100100","1111001001111010","1111001011010111","1111001100000110","1111000110101110","1111000000000000","1110111111111001","1111000101010111","1111001000011000","1111000101111010","1111000011100111","1111000111011100","1111010000111000","1111011011101000","1111100101001011","1111101101100100","1111110100101010","1111111001101001","1111111101100101","0000000100010111","0000010000100001","0000011110011000","0000100110111011","0000101000100001","0000101001011100","0000101111011100","0000111000001010","0000111101001101","0000111100110010","0000111010010110","0000111000111001","0000111000111011","0000111010001101","0000111011100101","0000111010010111","0000110101010011","0000101110101001","0000101000011001","0000100001101100","0000011010011100","0000010101000100","0000010001001001","0000001001011111","1111111101000000","1111110011000110","1111110000001010","1111101011110110","1111011101001110","1111001011001100","1111000100001101","1111000111111101","1111001000001001","1110111111111101","1110111011010000","1111000001011011","1111001000010010","1111000101000111","1110111110101111","1111000010000110","1111001101100101","1111010101000000","1111010101101001","1111011000101011","1111100010100001","1111101100011111","1111110001100011","1111110111000101","0000000011011011","0000010011010110","0000011110010001","0000100001011010","0000100001101000","0000100100100101","0000101011011111","0000110011111110","0000111010110010","0000111110001001","0000111110111011","0000111111010010","0000111111111011","0000111111011011","0000111101000000","0000111010001000","0000111000010000","0000110101111100","0000110000010010","0000100110111000","0000011101001011","0000010110110001","0000010011011001","0000001111010001","0000000111101010","1111111101100000","1111110011011011","1111101010110001","1111100011010101","1111011100101101","1111010110010001","1111001111000111","1111000111101100","1111000010011010","1111000000110100","1111000001010111","1111000001110001","1111000010010000","1111000100001000","1111000110110001","1111001000111011","1111001011100101","1111010000100001","1111010111000111","1111011101101011","1111100100010010","1111101011011011","1111110001111110","1111110111111001","0000000000001011","0000001011011101","0000010100100100","0000010111101000","0000011001100000","0000100001001001","0000101100100101","0000110100010000","0000110111011101","0000111011111101","0001000010010110","0001000100110100","0001000010000110","0000111111111010","0000111111111110","0000111100011101","0000110011000011","0000101010101101","0000101001011100","0000101011011111","0000101001100010","0000100001110111","0000010111000100","0000001011000110","1111111111101011","1111110110111010","1111110000001010","1111101000100000","1111100000100111","1111011100011101","1111011010111100","1111010101001011","1111001001110000","1111000001010101","1111000010010100","1111000110101100","1111000101010101","1110111111111101","1110111110111101","1111000011010110","1111000110101010","1111000111101010","1111001101001110","1111011010001100","1111100111000000","1111101100001110","1111101101110110","1111110101100101","0000000100010110","0000010000101111","0000010100100110","0000010110000001","0000011110010001","0000101011101100","0000110011101010","0000110010000001","0000101111011001","0000110100100000","0000111101101110","0001000001001011","0000111101010011","0000111001011100","0000111001100100","0000111001111101","0000111000010010","0000110111111011","0000111001101010","0000110111000000","0000101011101010","0000011101110010","0000010101101011","0000010001111101","0000001011100011","0000000001110111","1111111001111100","1111110011100001","1111101000111010","1111011010100111","1111010001001111","1111010000101101","1111010010000101","1111001110010110","1111001000010110","1111000110010001","1111000111101100","1111001000010010","1111000111010110","1111000110111111","1111000111010001","1111001000001100","1111001100100000","1111010101010001","1111011101111001","1111100010100010","1111100110101011","1111101111001001","1111111001000110","1111111110100100","0000000001011100","0000001001010111","0000010111010101","0000100011011011","0000101000000111","0000101000111101","0000101100000101","0000110010011111","0000111001010011","0000111110100110","0001000010000011","0001000010111011","0001000000100011","0000111100001011","0000111000110100","0000111000001010","0000110111101000","0000110010110011","0000101010000100","0000100011010000","0000100000101101","0000011011101110","0000001110010011","1111111110011100","1111110110101101","1111110101011011","1111101110111001","1111100000011010","1111010100101101","1111010010101100","1111010011111101","1111010000110001","1111001010001001","1111000011000010","1110111010110000","1110110011101011","1110110100101011","1110111101100000","1111000100100110","1111000101101000","1111000110111100","1111001011100101","1111001101100110","1111001101010100","1111010110001001","1111101010001011","1111111001001100","1111111000011010","1111110100111101","1111111111100101","0000010010110111","0000011110010011","0000100000001000","0000100010110000","0000101001010111","0000110000000111","0000111000010111","0001000011100010","0001001000010101","0000111110101100","0000110001011111","0000110010011000","0000111111010000","0001000100111111","0000111011100101","0000101110111110","0000101010011101","0000101010101110","0000100111011011","0000011110101111","0000010011111010","0000001010011110","0000000100110010","0000000001010011","1111111001111111","1111101100101010","1111100000100101","1111011100010000","1111011010011001","1111010010011110","1111000111110010","1111000100011100","1111000111111100","1111000111011101","1110111111100000","1110111001000010","1110111010111011","1111000001001001","1111000101011011","1111001000001000","1111001100001110","1111010001011111","1111010110111000","1111011101110101","1111100111101000","1111110010110010","1111111101010001","0000000110101010","0000001110110100","0000010101001111","0000011010011101","0000011111110010","0000100101101010","0000101100000001","0000110011100001","0000111011100101","0001000000101100","0000111111111111","0000111011111111","0000111010011010","0000111101010000","0001000000110111","0001000000110111","0000111100110001","0000110111000101","0000110001110111","0000101100110000","0000100101101010","0000011011110001","0000010001010000","0000001000101101","0000000001101000","1111111001110010","1111110001010110","1111101010000001","1111100010101001","1111011000101110","1111001110110101","1111001011000011","1111001101000011","1111001100101010","1111000101101000","1110111110011111","1110111110001010","1111000001010100","1111000000101111","1110111101101010","1110111111010000","1111000110111101","1111001111001100","1111010100110010","1111011001111111","1111100000010100","1111100110010101","1111101100011101","1111110101101111","0000000010001110","0000001101010100","0000010011111101","0000011000100000","0000011110110010","0000100110111010","0000101110001110","0000110011100001","0000111000000100","0000111100111011","0001000000101001","0001000001000101","0000111111000111","0000111110001000","0000111110100111","0000111100000011","0000110011101111","0000101010100101","0000100110111110","0000100110111010","0000100010111101","0000011001110011","0000010001001111","0000001011011011","0000000011110001","1111111000110000","1111101111101101","1111101010111111","1111100101000011","1111011010011010","1111010001000010","1111001111010001","1111010001101101","1111010001001001","1111001101010010","1111001010001010","1111000111100101","1111000011010000","1110111111111010","1111000001111111","1111000111001101","1111001001011110","1111001001101100","1111001111010001","1111011011111010","1111100111100101","1111101011110100","1111101100111100","1111110011100000","0000000000101001","0000001101110100","0000010110001000","0000011011010101","0000100001101011","0000101010101001","0000110100101111","0000111101011011","0001000010011010","0001000010110000","0001000000011000","0000111110100110","0000111110011011","0000111101100001","0000111010001010","0000110110000101","0000110011010111","0000110001000001","0000101100111011","0000100111010110","0000100001001111","0000011001000001","0000001101010111","0000000001101101","1111111011011001","1111111010000101","1111110111101111","1111110000101101","1111100111101101","1111100000100011","1111011011000001","1111010100110010","1111001101010000","1111000101110100","1111000000100000","1110111111011010","1111000010010100","1111000100101001","1111000001101110","1110111100000001","1110111011100001","1111000011001100","1111001101011000","1111010100101011","1111011010111110","1111100011110001","1111101101000001","1111110011010100","1111111000111000","0000000010000100","0000001101001001","0000010100110011","0000011000111000","0000011110010011","0000100110101010","0000101110100011","0000110100000100","0000111000100111","0000111011101100","0000111010111101","0000111000100001","0000111010000011","0000111111001101","0001000000010000","0000111001011101","0000110001001010","0000101101101111","0000101100001000","0000100110010100","0000011101100000","0000010110100110","0000010001000010","0000001001000110","0000000000011001","1111111011001011","1111110110110011","1111101100010100","1111011100110100","1111010001101111","1111001111000001","1111001101101100","1111000111110010","1111000001001110","1110111111100000","1111000000010111","1110111111100011","1110111111110111","1111000101110001","1111001101010010","1111001111001010","1111001110000111","1111010011111110","1111100001001110","1111101010101001","1111101011000000","1111101100001001","1111110111010110","0000000110000010","0000001100001101","0000001011101111","0000010001000111","0000011110111011","0000101010000100","0000101011100101","0000101011000011","0000110001100000","0000111011111001","0001000001100001","0001000001101000","0001000010000001","0001000100001010","0001000011100000","0000111101111111","0000110111001111","0000110010101100","0000101111001010","0000101001111000","0000100010100001","0000011010011001","0000010010011001","0000001010110111","0000000100001101","1111111110000100","1111110110100101","1111101100000001","1111011111100111","1111010101101111","1111010001011110","1111010000010010","1111001100100000","1111000100101011","1110111101100100","1110111011101001","1110111101100110","1111000000000011","1111000010100010","1111000101001111","1111000101110101","1111000011110110","1111000100100010","1111001100001101","1111010110101101","1111011101110010","1111100011011010","1111101101100001","1111111001111000","0000000000110011","0000000011010001","0000001010110110","0000011001100100","0000100101100111","0000101000101011","0000101001000111","0000101110010010","0000110101010100","0000111000010101","0000111001001111","0000111101010100","0001000011011111","0001000101111101","0001000010000010","0000111001111011","0000110001011011","0000101100101111","0000101110000010","0000110001001010","0000101101011111","0000100000000000","0000001111110010","0000000101110010","0000000011010110","0000000010111101","1111111110100111","1111110011110111","1111100101011001","1111011010001000","1111010110111000","1111011000001000","1111010110010001","1111001111011010","1111000111110110","1111000010000110","1110111101001110","1110111010110111","1110111110110011","1111000111011000","1111001110000010","1111010001000101","1111010101010101","1111011100011101","1111100001100100","1111100010011000","1111100011111101","1111101010110011","1111110100011010","1111111100110100","0000000100100011","0000001101101011","0000010111110011","0000100001101001","0000101010011111","0000110000000100","0000110000001111","0000101110100000","0000110001110110","0000111010110010","0001000001110011","0001000010001111","0001000000011001","0001000000111110","0001000001000011","0000111100001001","0000110100010110","0000101110011001","0000101001011101","0000100001110101","0000011000111011","0000010011001001","0000001111001101","0000000111001110","1111111010111000","1111110001011001","1111101110110111","1111101101100111","1111100110100100","1111011011011101","1111010011011111","1111010000110000","1111001110010001","1111001000010010","1111000001011110","1110111110101011","1111000000101111","1111000100001100","1111000101110100","1111000110010010","1111001001110001","1111010010111111","1111011110111110","1111100111001101","1111101001010101","1111101010001111","1111101111101001","1111111001000110","0000000010011000","0000001010010100","0000010010110001","0000011011011000","0000100001100110","0000100110000000","0000101100101100","0000110110101001","0000111110111000","0001000000001011","0000111011101100","0000110111110101","0000111001110111","0001000000011110","0001000100011000","0000111111000110","0000110010100010","0000101000001001","0000100110011011","0000101001000101","0000100110111001","0000011101010110","0000010001111111","0000001001011100","0000000010100010","1111111010100111","1111110010000110","1111101010101010","1111100100010101","1111011110001111","1111010111110100","1111010000011111","1111001000010100","1111000001100101","1110111111000010","1111000000001010","1111000001111010","1111000011000111","1111000100110111","1111000110101101","1111000110011110","1111000101010000","1111000111110000","1111010000000100","1111011010100110","1111100011100101","1111101011100001","1111110011111111","1111111100001110","0000000011111010","0000001101000000","0000010111010000","0000011110011110","0000100001010101","0000100100110111","0000101100100010","0000110011101101","0000110101011000","0000110101001000","0000111000110010","0000111101101000","0000111101000001","0000111000100101","0000110111110000","0000111010110100","0000111010011010","0000110011110011","0000101011100001","0000100100010000","0000011100010001","0000010100100010","0000010000001011","0000001100001111","0000000010010110","1111110100100101","1111101011111010","1111101001011011","1111100100011110","1111011010000001","1111010001111111","1111010000101101","1111001111000101","1111000111001111","1110111110110100","1110111100110011","1110111110001100","1110111100110100","1110111010111001","1110111111010111","1111001010101110","1111010110011011","1111011101000100","1111011110100111","1111011110110000","1111100001111110","1111101001111101","1111110011101001","1111111011011111","0000000010110001","0000001100100001","0000010110011010","0000011011100101","0000011101111110","0000100100110110","0000110000110111","0000111001011111","0000111001001001","0000110101010110","0000110110110110","0000111110100000","0001000101000110","0001000011111100","0000111011010100","0000110010001000","0000101110011101","0000101101111101","0000101000100111","0000011101001110","0000010100110100","0000010101000001","0000010101100011","0000001011111010","1111111011110010","1111110001000111","1111101101011001","1111100111011010","1111011100001001","1111010011001101","1111010000101100","1111001110110001","1111001001001111","1111000100110011","1111000101010010","1111000101111101","1111000001111010","1110111101001110","1110111110001111","1111000011011000","1111000110111000","1111001000110001","1111001110000010","1111010111100001","1111100000101110","1111100111010101","1111101101110010","1111110101100111","1111111100111000","0000000011010001","0000001100011011","0000011001101100","0000100101010001","0000101000110111","0000100111100100","0000101010110101","0000110101100101","0001000000001100","0001000011101100","0001000010110110","0001000011101000","0001000101010001","0001000011000101","0000111101101100","0000111001101111","0000110110110001","0000101111110010","0000100101000100","0000011101010001","0000011010100100","0000010110100001","0000001100101010","0000000010010001","1111111101101101","1111111011110101","1111110100110100","1111100111111111","1111011011110101","1111010011110100","1111001101100110","1111001000001111","1111000110110100","1111001001100001","1111001010001111","1111000100010101","1110111100010011","1110111010010110","1110111111011000","1111000100010101","1111000100110110","1111000101010101","1111001011111101","1111010111011000","1111100000101011","1111100101010010","1111101010010001","1111110100101110","0000000010100011","0000001101001101","0000010010000101","0000010101010100","0000011100000101","0000100101110100","0000101101000110","0000101111000111","0000110000000101","0000110101111001","0000111110111111","0001000010111010","0000111101101110","0000110101111111","0000110011111100","0000110110010000","0000110101011101","0000110000001101","0000101100100001","0000101100110110","0000101011100000","0000100011100001","0000010111101100","0000001101010011","0000000100101110","1111111011100011","1111110001111100","1111101001100001","1111100001110000","1111011001101100","1111010011000011","1111001111110101","1111001101111010","1111001000110010","1111000000000010","1110111001000101","1110111001001000","1110111110101111","1111000011010110","1111000011100000","1111000011100111","1111001001100010","1111010011001000","1111011000101110","1111011010000011","1111100000011110","1111101111111001","1111111101101011","1111111111010001","1111111011101011","0000000010011100","0000010100010001","0000100001111001","0000100010110111","0000100000011101","0000100101101100","0000110000000011","0000110110111100","0000111001101101","0000111101110010","0001000011111111","0001000111001111","0001000011110010","0000111011000110","0000110010000101","0000101101110100","0000101111001100","0000110000001010","0000101001110000","0000011101111110","0000010110000001","0000010100110000","0000010010000111","0000000111110111","1111111011001001","1111110011001111","1111101101100011","1111100011000111","1111010101000110","1111001010111010","1111000110100100","1111000011011011","1110111111110001","1110111110111010","1111000001101000","1111000011101100","1111000010100101","1111000000101011","1111000000011010","1111000001101010","1111000100110111","1111001011010010","1111010011010101","1111011001110100","1111011111100111","1111101000011011","1111110011001001","1111111010010001","1111111101011010","0000000011010110","0000001111011001","0000011011100011","0000100001101001","0000100100000110","0000101000101010","0000101111100101","0000110101100101","0000111010000011","0000111101111100","0001000000000110","0000111111100100","0000111110001001","0000111100011010","0000110111100010","0000101111100110","0000101010100100","0000101011000111","0000101010001000","0000100000100110","0000010010111110","0000001010100000","0000000111000101","0000000001100110","1111111000110111","1111110001110000","1111101011111101","1111100010000001","1111010100111001","1111001100010011","1111001001100000","1111000100111000","1110111100000101","1110110111101110","1110111100111100","1111000011110100","1111000011110010","1111000001001111","1111000101001010","1111001101011010","1111010000101011","1111001110100010","1111010000100000","1111011011011000","1111101001001111","1111110011010000","1111111001011100","1111111110101011","0000000011110100","0000001001101000","0000010001111101","0000011011110011","0000100011001111","0000100111010010","0000101011011001","0000110001001010","0000110101101000","0000110111100101","0000111010100100","0001000000001011","0001000011100011","0001000000110011","0000111100000111","0000111011101010","0000111101011000","0000111001101000","0000101110110101","0000100011110111","0000011110001100","0000011010111000","0000010011101101","0000000111100011","1111111010110101","1111110001100101","1111101011110001","1111100111001111","1111100011000000","1111011110101111","1111011000100110","1111001110101101","1111000011100011","1110111101010101","1110111110011101","1111000001101100","1111000001010101","1110111111001001","1111000000010010","1111000100010001","1111000110101110","1111001000100010","1111001111000011","1111011001111100","1111100010001001","1111100101001100","1111101001100001","1111110011110011","1111111111001111","0000000101110111","0000001010010011","0000010010011100","0000011101001100","0000100100110000","0000101000001111","0000101011111000","0000110000101101","0000110011100110","0000110100101100","0000111000101000","0001000000100001","0001000110011001","0001000101010101","0001000000001100","0000111100010101","0000111001000001","0000110001100000","0000100101101111","0000011011110110","0000010111111011","0000010111000010","0000010011101011","0000001100001100","0000000010101011","1111111001000100","1111101111110111","1111100111001111","1111011111010011","1111011000001101","1111010010111000","1111010000011100","1111001111111100","1111001110010111","1111001010001100","1111000101100111","1111000011001010","1111000010011100","1111000010001101","1111000100001000","1111001010100101","1111010011001111","1111011000000001","1111010111011010","1111010111111101","1111100000011011","1111101110011000","1111111001001100","1111111110001110","0000000100001110","0000010000100101","0000011110101101","0000100110101010","0000101000101010","0000101011000100","0000101111011101","0000110001101011","0000110001011110","0000110100010110","0000111100000101","0001000010011101","0001000010000110","0000111100111011","0000110111100001","0000110011101110","0000110010101111","0000110101000000","0000110101101010","0000101101100010","0000011110010101","0000010010100011","0000001110000000","0000001000001100","1111111011001100","1111101110010111","1111101001110010","1111101000100110","1111100001011011","1111010101010010","1111001011110100","1111000110111110","1111000011111000","1111000010111010","1111000101010101","1111000111011101","1111000110001100","1111000101100101","1111001001001111","1111001100010011","1111001010011000","1111001010000011","1111010010110100","1111011110011100","1111100001101010","1111011111101101","1111100110001011","1111110110101001","0000000011100011","0000000101100011","0000000101111010","0000001110110011","0000011100101011","0000100110011011","0000101011010110","0000110001001001","0000111001001000","0000111110101101","0000111111001000","0000111101100011","0000111110111100","0001000011010110","0001000100101111","0000111101101010","0000110001011011","0000101001101111","0000101010010011","0000101011010101","0000100100101001","0000011001011000","0000010001111110","0000001110011111","0000000111100110","1111111011100101","1111110001000110","1111101100000110","1111101000000001","1111100000000001","1111010110010101","1111001111110111","1111001100101110","1111001000110100","1111000001111001","1110111010110111","1110111001011000","1110111111010000","1111000110001100","1111000101111001","1111000000000111","1111000000010101","1111001011111111","1111011001101100","1111011111011000","1111100001011001","1111101001110110","1111110111000110","1111111111011100","0000000010010010","0000001000000010","0000010010000101","0000011001000110","0000011011101100","0000100001100111","0000101101010110","0000110111010110","0000111010110100","0000111100011001","0001000000000111","0001000011011000","0001000100000010","0001000011111000","0001000010000100","0000111011010011","0000110010011110","0000101110101100","0000101110010110","0000101000010001","0000011100100110","0000010110011011","0000010111111111","0000010011111111","0000000010101001","1111101111100010","1111100111110010","1111100110011010","1111011111010010","1111010011111011","1111001110111010","1111010000101101","1111001111011101","1111001000010000","1111000011000000","1111000100001101","1111000101101111","1111000001100011","1110111011100110","1110111100100101","1111000110000100","1111010000011110","1111010011111110","1111010001111010","1111010011010011","1111011101101111","1111101100000000","1111110101001111","1111111001001100","1111111111001101","0000001001110001","0000010010111110","0000010111101111","0000011101101111","0000101001011111","0000110101111001","0000111011111110","0000111101000000","0000111101110011","0000111101110011","0000111010110000","0000111000110011","0000111100110101","0001000010001001","0001000000000001","0000111000000110","0000110100000001","0000110100101010","0000101111111110","0000100001111010","0000010100001100","0000001111010110","0000001110010101","0000001000000000","1111111101000101","1111110100010010","1111101110011111","1111100111001110","1111011101011011","1111010100001000","1111001100100101","1111000110000011","1111000001101001","1111000000100110","1111000000101110","1110111111001100","1110111101011101","1110111111000000","1111000011101010","1111001000010001","1111001011011101","1111001110101001","1111010011101000","1111011011011101","1111100101111001","1111110000010011","1111110111100100","1111111100001110","0000000001101111","0000001001000111","0000010000011010","0000010111110101","0000100001100111","0000101100010110","0000110011101011","0000110111110010","0000111100111110","0001000010011011","0001000001111000","0000111011001101","0000110111010010","0000111010111111","0000111111110000","0000111101111011","0000110110111011","0000101111110110","0000101001010101","0000100010100010","0000011101001100","0000011000110001","0000010000011110","0000000011110110","1111111010011000","1111111000100100","1111110111111110","1111110000110011","1111100101001100","1111011100010001","1111010111010011","1111010010101110","1111001100111100","1111000110011001","1110111111010010","1110111010000111","1110111011010101","1111000001110001","1111000101100101","1111000011011101","1111000001101100","1111000101011011","1111001010110111","1111001110100101","1111010101101001","1111100011101110","1111110001100001","1111110111010101","1111111010100110","0000000101011011","0000010101110000","0000100000011001","0000100010010010","0000100011010100","0000101001001010","0000110001010100","0000111000010001","0000111101110101","0001000001111101","0001000011111011","0001000100111011","0001000101100101","0001000010100110","0000111001101110","0000110000001010","0000101100110010","0000101101111101","0000101100000001","0000100100101011","0000011100110001","0000010111101000","0000010011010110","0000001101001000","0000000100000110","1111111000011010","1111101100011111","1111100100101111","1111100001100011","1111011100111011","1111010011010010","1111001001110111","1111000101111110","1111000011110000","1110111110011100","1110111011100100","1111000010010010","1111001100010000","1111001100100110","1111000100001100","1111000000110101","1111001000010001","1111010001101111","1111010110101011","1111011011110011","1111100101100000","1111101111100110","1111110110010001","1111111101000001","0000000110101100","0000010000000100","0000010111000011","0000011111000011","0000101000111101","0000101111011010","0000110000011000","0000110010000101","0000111000111001","0001000000010011","0001000011010111","0001000100011000","0001000110011001","0001000110100011","0001000010101011","0000111110110101","0000111101101110","0000111010000101","0000101111010011","0000100010100011","0000011011000100","0000010111000100","0000010000001011","0000000110001100","1111111101000010","1111110100010001","1111101001011011","1111011111100001","1111011010111111","1111011000101101","1111010010000000","1111001000100010","1111000100011000","1111000110011100","1111000110100001","1111000001000000","1110111101000110","1111000001000011","1111001000000010","1111001010000000","1111001000000011","1111001010000101","1111010010110111","1111011101001001","1111100011111111","1111101000010010","1111101101011101","1111110101000110","1111111111000011","0000001010100001","0000010101010100","0000011101000000","0000100001111010","0000100111000111","0000101110000010","0000110100010100","0000110111011100","0000111000010010","0000111001011100","0000111100000011","0000111111111100","0001000100001110","0001000110000010","0001000001110010","0000111000010101","0000110000001101","0000101110000001","0000101110000110","0000101001100101","0000011111101011","0000010101010100","0000001101011001","0000000110000101","1111111101100100","1111110100101101","1111101100110010","1111100101110010","1111011111100001","1111011001101111","1111010011101111","1111001101101000","1111001000110011","1111000101100001","1111000010000110","1110111111000010","1111000000010101","1111000111000110","1111001101000100","1111001100010001","1111001000001001","1111001001000111","1111010000101001","1111011000011001","1111011101000001","1111100010110001","1111101101111011","1111111011110000","0000000101110111","0000001001111001","0000001011101110","0000010001011011","0000011101001100","0000101010011100","0000110010001110","0000110011100000","0000110100100011","0000111010000001","0001000000010101","0001000001101010","0000111110111111","0000111101101111","0000111110010101","0000111011100101","0000110011100000","0000101010111110","0000100111000011","0000100110110001","0000100101001010","0000011111001011","0000010101111100","0000001100100100","0000000100011011","1111111011111100","1111110001011011","1111100110111100","1111100000010011","1111011101010011","1111011001001011","1111010001110001","1111001010111001","1111000111101100","1111000101000100","1110111111001110","1110111001100110","1110111010011111","1111000000101011","1111000100011010","1111000011001010","1111000011111110","1111001100111011","1111011001110111","1111100001110100","1111100011001010","1111100101100010","1111101111100100","1111111110011011","0000001001110110","0000001110100000","0000010001000010","0000010110101100","0000011110101001","0000100101010101","0000101011001001","0000110010111010","0000111010110101","0000111101010011","0000111001111010","0000110111111100","0000111100000100","0001000000111010","0000111110101001","0000110110010111","0000101111101000","0000101101000000","0000101001111000","0000100011011001","0000011100101011","0000011000010101","0000010011011110","0000001010100000","1111111110111110","1111110100111011","1111101100110100","1111100100011101","1111011100001111","1111010111000111","1111010101001111","1111010010011010","1111001011101111","1111000100000111","1111000000100010","1111000001100010","1111000010111010","1111000010001101","1111000010001101","1111000110010101","1111001100011111","1111001111000001","1111001100111000","1111001100101111","1111010101010110","1111100100100111","1111110001110010","1111111000010011","1111111100010010","0000000011000011","0000001011100110","0000010010010100","0000011000001010","0000100000100001","0000101001011111","0000101101110000","0000101110010111","0000110011000111","0000111110001111","0001000111011111","0001001000000111","0001000100110011","0001000100111111","0001000110001011","0001000001011001","0000111000011010","0000110011001101","0000110001100011","0000101010110001","0000011100111000","0000010000111100","0000001100110000","0000001001110111","0000000000100001","1111110011011001","1111101010001011","1111100110001010","1111100010110010","1111011101101001","1111010111101010","1111010001001100","1111001010001111","1111000100101111","1111000010010101","1111000001110010","1111000001101011","1111000011001101","1111000111000100","1111001010110100","1111001100011101","1111001101111011","1111010001010101","1111010101011000","1111011001011011","1111100001000110","1111101110011101","1111111011110000","0000000010010010","0000000101000010","0000001100111111","0000011010110110","0000100101000110","0000100110010011","0000100101011110","0000101011001001","0000110100101101","0000111001000111","0000110111010010","0000110111101110","0000111111100111","0001001000100110","0001001000011011","0000111101110000","0000110001100001","0000101100000110","0000101100011001","0000101010110001","0000100010110001","0000010111100011","0000001110010100","0000000111101000","0000000000011110","1111111000010001","1111110010000011","1111101111001100","1111101100011101","1111100101101110","1111011010100101","1111001110001111","1111000100101110","1111000000100100","1111000000111001","1111000001011000","1110111110110001","1110111011101110","1110111101011001","1111000011010100","1111000111110110","1111001001101010","1111001110000111","1111010111011011","1111011111100011","1111100010001100","1111100101001000","1111101111000001","1111111011110000","0000000010111001","0000000101010101","0000001010100010","0000010011011010","0000011010100101","0000011111111110","0000101000100101","0000110010011111","0000110101011111","0000110001101111","0000110001110000","0000111001110001","0001000000100110","0000111111000110","0000111011101101","0000111110010011","0001000010000001","0000111101010001","0000110001011010","0000100111011010","0000100001010101","0000011001110111","0000001111111111","0000001000101011","0000000100101110","1111111110100101","1111110100001110","1111101010110000","1111100101101010","1111100001001001","1111011001000000","1111001111100000","1111001001000000","1111000101011000","1111000010000111","1110111111100100","1110111111100011","1111000000101110","1111000000010100","1110111111010110","1111000001001101","1111000101111111","1111001010100111","1111001110111011","1111010110100000","1111100010001011","1111101101000101","1111110011001001","1111110110101000","1111111100010010","0000000101000100","0000001110111101","0000011001011110","0000100100110100","0000101110010101","0000110010011111","0000110010011111","0000110011110001","0000111001000011","0000111110110001","0001000000011001","0000111110100010","0000111101100010","0000111111010010","0001000000011001","0000111100010001","0000110010100001","0000100111011010","0000011110110000","0000011000010101","0000010010000001","0000001011111111","0000001000001001","0000000101100010","1111111111111111","1111110101010100","1111101000110111","1111011111101110","1111011010101001","1111010101100100","1111001101000100","1111000011010001","1110111110000010","1111000000000101","1111000100110110","1111000101100111","1111000010100100","1111000010101000","1111001000110000","1111001110011111","1111001101100110","1111001010100001","1111001110001011","1111011000011110","1111100001000101","1111100101001001","1111101010101111","1111110101010100","1111111111100100","0000000100111100","0000001001001100","0000010000111110","0000011001100001","0000011110100011","0000100011000100","0000101100001011","0000110110111100","0000111011110110","0000111010110111","0000111011001011","0000111111000101","0001000000101001","0000111100110010","0000111001001001","0000111010011010","0000111011101001","0000110110000000","0000101011111010","0000100100110111","0000100001000110","0000011001011010","0000001011001110","1111111100101010","1111110011000011","1111101100101101","1111100110110101","1111100010101011","1111100000001010","1111011010000000","1111001101100101","1111000010000010","1111000000000010","1111000101000001","1111000110011011","1111000000011111","1110111010011001","1110111011011010","1111000010100111","1111001010110110","1111010000110100","1111010011100110","1111010100011110","1111010111110110","1111100001000000","1111101100000000","1111110001101001","1111110010100010","1111110111011100","0000000100000100","0000010001001000","0000010111110000","0000011011100000","0000100011001000","0000101101100110","0000110101001111","0000111001011111","0000111101010110","0000111111101101","0000111101011001","0000111001001100","0000111001000101","0000111011101100","0000111001001010","0000110000000011","0000101001000111","0000101010001010","0000101100101001","0000100110111100","0000011001111010","0000001110011101","0000001000010011","0000000010010110","1111111000001011","1111101100001110","1111100010110000","1111011100000111","1111010110110100","1111010011011010","1111010010000110","1111001111101010","1111001001001000","1111000001001101","1110111101101000","1110111111100100","1111000010110101","1111000100101110","1111000111010010","1111001100011010","1111010010010101","1111010110111011","1111011010110011","1111011110101110","1111100001111010","1111100101110111","1111101111010101","1111111111000010","0000001100101110","0000001111111011","0000001100011001","0000001110110010","0000011100011010","0000101100110000","0000110101100010","0000110111010110","0000111001100000","0000111110011011","0001000001111010","0001000001001111","0000111110101101","0000111100111110","0000111011101010","0000111001111111","0000111000011111","0000110110101001","0000110001110110","0000101000100001","0000011100011101","0000010000110010","0000000111011000","0000000000111101","1111111100100110","1111110110100101","1111101011100100","1111011110010100","1111010110100100","1111010110111110","1111011000000110","1111010001101011","1111000101111111","1110111111001101","1111000010000101","1111001000000111","1111000111110011","1110111111010111","1110110110000111","1110110101000100","1110111110101101","1111001101000001","1111010111100010","1111011011100001","1111011101011111","1111100010110010","1111101011111100","1111110101110101","1111111110001011","0000000101000001","0000001011101101","0000010011101001","0000011100100101","0000100100001000","0000101000111011","0000101101011111","0000110100100011","0000111011101111","0000111110101010","0000111110110010","0001000001101000","0001000110110001","0001000111010110","0001000001011101","0000111011011110","0000111000110110","0000110100011110","0000101010110111","0000100001011011","0000011100101010","0000010111101101","0000001101010110","0000000010001011","1111111100011110","1111111000100110","1111101111100110","1111100100001000","1111011101011010","1111011001111000","1111010010110111","1111001010011101","1111001000010101","1111001010011100","1111000110011101","1110111011110111","1110110110101110","1110111101001000","1111000110001011","1111001000111010","1111001001001000","1111001110001100","1111010110100101","1111011100111100","1111100001110110","1111101000010101","1111101110010101","1111110001010110","1111110110010100","0000000011100010","0000010100111100","0000011111100101","0000100000101011","0000100001001110","0000101000100111","0000110011000010","0000111000101111","0000111001000110","0000111001100111","0000111100111011","0001000000001100","0001000000101100","0000111111001001","0000111100111010","0000111001111100","0000110110100010","0000110011101010","0000101111111010","0000100111100101","0000011010011001","0000001101110110","0000000110011001","0000000001100000","1111111010000110","1111110000100110","1111101001010001","1111100100010110","1111011101101001","1111010011110110","1111001010110110","1111000101111110","1111000100011001","1111000100000010","1111000100001000","1111000100001001","1111000011101001","1111000011101001","1111000101001001","1111000111000101","1111001001001010","1111001110011100","1111011000011011","1111100001110111","1111100101000111","1111100101101001","1111101011100111","1111110110111101","1111111111110010","0000000100011001","0000001100101010","0000011100001011","0000101010101110","0000110000001000","0000101111101110","0000110001110000","0000110111011001","0000111100001010","0000111110000101","0000111110001000","0000111100011000","0000111010000101","0000111011100011","0001000001011001","0001000011111100","0000111100010000","0000101111001001","0000100110111101","0000100100101100","0000011111110001","0000010100010001","0000001000001111","0000000000111001","1111111011010001","1111110011010101","1111101011001011","1111100101110111","1111100000101100","1111011000000010","1111001110101000","1111001001010111","1111000110111001","1111000010001101","1110111100000000","1110111010010001","1110111110011001","1111000010101011","1111000011010100","1111000100000000","1111001001000101","1111010000010000","1111010100100111","1111010110100001","1111011011000101","1111100100100110","1111101111110010","1111111000011011","1111111101111110","0000000011001101","0000001010111110","0000010101101001","0000100000100100","0000101000010001","0000101011101101","0000101101011100","0000110000111001","0000110111001001","0000111110010110","0001000011001111","0001000011010010","0000111111000101","0000111011001110","0000111100010011","0001000000100000","0001000000000000","0000110101111110","0000100111010101","0000011101001011","0000011001111000","0000010111010111","0000010000000000","0000000100101000","1111111001001110","1111101111011110","1111100111001111","1111100001000100","1111011100110011","1111010111101010","1111001111000101","1111000101000110","1110111110110101","1110111110110000","1111000010001100","1111000100101011","1111000100001000","1111000001110111","1111000001000111","1111000100001011","1111001010000110","1111001111100011","1111010010111101","1111010110011111","1111011101000001","1111100110111000","1111110010101010","1111111111000011","0000001001011010","0000001110000111","0000001110000010","0000010000101111","0000011011111101","0000101010110100","0000110011010100","0000110011101000","0000110011011101","0000111000000011","0000111101111001","0001000000001011","0001000000000000","0001000000101000","0001000001100101","0001000000001101","0000111011101100","0000110100011100","0000101010101010","0000100000001100","0000011000100010","0000010100011011","0000010000001111","0000001000110111","1111111111101110","1111110111100001","1111110000011011","1111101001010111","1111100010000100","1111011001111100","1111010000010010","1111000111101111","1111000101001000","1111001000000100","1111001001011010","1111000100101010","1110111110011100","1110111101010001","1111000000001100","1111000010001000","1111000011000100","1111000111001110","1111001111010001","1111010111100111","1111011110011000","1111100100110000","1111101011001101","1111110001101010","1111111010000001","0000000101100101","0000010001000010","0000011000011011","0000011101101001","0000100101001010","0000101101101010","0000110001111110","0000110010100101","0000110101101011","0000111100111111","0001000010111001","0001000011001111","0001000000001111","0000111101000100","0000111001111000","0000110110111110","0000110101010001","0000110010011101","0000101011010111","0000100010111110","0000011111001010","0000011101010111","0000010100011001","0000000011101101","1111110101111001","1111110000001101","1111101011011001","1111100010011111","1111011100001001","1111011100011000","1111011001110001","1111001101000111","1111000000110111","1111000010000011","1111001010010001","1111001001110001","1111000001100011","1111000000101110","1111001010000100","1111001111110101","1111001011110101","1111001001011011","1111010001111000","1111011110110011","1111100111101000","1111101110110010","1111111000010100","1111111111011101","1111111111111000","0000000000001101","0000001000101010","0000010101101111","0000011110001001","0000100001000011","0000100101100011","0000101110111101","0000111001101011","0001000001100111","0001000101000110","0001000011110100","0001000000000100","0000111110110010","0001000001000110","0001000001010000","0000111010101110","0000110001111100","0000101101110010","0000101100101010","0000100111000110","0000011011100101","0000010000111100","0000001100010101","0000001010011101","0000000100100011","1111111000100101","1111101011000100","1111100001111101","1111011110100111","1111011100101101","1111010111100100","1111001111110101","1111001001100100","1111000101111101","1111000011000100","1111000000111100","1111000001010001","1111000010001001","1111000000000110","1110111110010000","1111000100010111","1111010010010011","1111011110001101","1111100010110011","1111100110000010","1111101100100011","1111110001010110","1111110001011101","1111110101000101","0000000010011001","0000010000100110","0000010101001110","0000010110001111","0000100000000111","0000101111111001","0000111000001101","0000111000001010","0000111011001010","0001000010101110","0001000011111000","0000111100110010","0000111001101011","0000111110101101","0000111111110011","0000110110110011","0000101111101110","0000110011101100","0000110111111011","0000101111110011","0000100001100000","0000011000110000","0000010001010110","0000000001000111","1111101110000011","1111100110100100","1111101000111100","1111100110010111","1111011100000010","1111010101110101","1111010111010011","1111010101000110","1111001001100010","1110111110110101","1110111110010111","1111000011001001","1111000100100001","1111000011001111","1111000100001000","1111000110110001","1111001000110001","1111001011110101","1111010010000011","1111011001011100","1111011111111111","1111100111001010","1111101111110010","1111110111100101","1111111110001000","0000000110101101","0000010010000011","0000011011110000","0000100001010001","0000100110001011","0000101101100101","0000110100001111","0000110101110100","0000110100001000","0000110100111111","0000111010101010","0001000001101101","0001000100110001","0001000001001110","0000111001011101","0000110011001011","0000110001000000","0000101110101101","0000100110110000","0000011010101011","0000010001010000","0000001100101100","0000001000001010","1111111111110110","1111110110011010","1111110000001000","1111101100110100","1111101000111001","1111100010001000","1111011001001011","1111010000100001","1111001010101100","1111000111110100","1111000101000111","1111000000101100","1110111100111100","1110111101011000","1111000001010111","1111000101100100","1111001001001000","1111001101011110","1111010001111110","1111010100111000","1111010111111011","1111011110011010","1111100111001111","1111101110101111","1111110110001101","0000000010001000","0000010000000111","0000010111011101","0000010110110111","0000011000011001","0000100010010100","0000101100111010","0000101111010000","0000101110100000","0000110101011001","0001000001111011","0001001000000111","0001000100100011","0000111111110001","0000111110110010","0000111100101010","0000110110001001","0000110000000100","0000101101100011","0000101001101001","0000100000100010","0000010111001001","0000010011000101","0000010001100001","0000001100001001","0000000010001111","1111110111011001","1111101101110100","1111100101111011","1111011111110010","1111011001001001","1111001111010001","1111000100111000","1111000000101110","1111000011011011","1111000101110010","1111000011110010","1111000010000000","1111000100000101","1111000110111110","1111001000111000","1111001110001101","1111011000001101","1111011111101010","1111100000001111","1111100001000100","1111101001110011","1111110110100110","1111111111001111","0000000100000011","0000001010110000","0000010100000011","0000011100110100","0000100100111101","0000101101001101","0000110010101110","0000110100001100","0000110110100111","0000111101110101","0001000100101011","0001000100011011","0000111111010111","0000111100100100","0000111100111010","0000111011110001","0000110111011110","0000110001100011","0000101010000110","0000100001100110","0000011100000011","0000011011011101","0000011010010100","0000010010000100","0000000100100000","1111111000101010","1111110000100011","1111101000101111","1111011111101011","1111010111100011","1111010001101110","1111001101011101","1111001010100001","1111001000101101","1111000110001100","1111000001111110","1110111110011011","1110111110010011","1111000000101100","1111000010111111","1111000100011010","1111000101101000","1111000111101000","1111001101001001","1111011000111111","1111101000010011","1111110011001000","1111110110100001","1111111000111111","0000000000111100","0000001011100111","0000010011010010","0000011001001110","0000100010010111","0000101101110011","0000110110001001","0000111010001111","0000111101001101","0000111111100100","0000111111110100","0001000000011100","0001000101000110","0001001010000000","0001000110100010","0000111010001000","0000101110111010","0000101100001110","0000101101010101","0000101001001110","0000011110110010","0000010100001101","0000001101010000","0000000111100001","1111111111110000","1111110110111011","1111110000001010","1111101011001001","1111100011010011","1111010110010010","1111001001010000","1111000011101011","1111000100110100","1111000100000101","1110111101011011","1110110111110110","1110111011000100","1111000100010010","1111001010100110","1111001010101110","1111001000100000","1111001000001110","1111001100000110","1111010101010111","1111100001101100","1111101010100010","1111101101010010","1111110000010110","1111111010000101","0000000110110010","0000001111000001","0000010011111010","0000011011101111","0000100101100011","0000101010110100","0000101100000110","0000110001001111","0000111011111010","0001000011111100","0001000011101011","0000111111010110","0000111101010111","0000111110010110","0000111111000001","0000111100110010","0000110110010010","0000101100101011","0000100101001100","0000100011110010","0000100100010011","0000011110101101","0000010010010000","0000000101101110","1111111100101111","1111110100000100","1111101001100111","1111100000101011","1111011011011001","1111010110011101","1111001111000100","1111001000001000","1111000101100111","1111000110001100","1111000101000010","1111000000010100","1110111010111111","1110111001100000","1110111101111110","1111000110011110","1111001110100100","1111010011001001","1111010101001011","1111011000100010","1111100000011010","1111101100111010","1111111010100000","0000000011110100","0000000110100111","0000000111100110","0000001101110011","0000011001110000","0000100100111011","0000101011001000","0000101111011000","0000110101001101","0000111010011110","0000111011101100","0000111010010111","0000111010110010","0000111110010100","0001000011001110","0001000111000100","0001000110101110","0000111111100011","0000110011110111","0000101010011111","0000100110111100","0000100101100111","0000100001101101","0000011010100111","0000010000111101","0000000100010100","1111110111001000","1111101111000011","1111101100011010","1111100111001010","1111011010001000","1111001100000100","1111000111000010","1111001010101111","1111001110001001","1111001011011111","1111000100100111","1110111110000010","1110111011011101","1110111110110010","1111000101100110","1111001010000011","1111001010011110","1111001100010101","1111010011100011","1111011011101000","1111011111100001","1111100011000011","1111101100111001","1111111010111010","0000000101010000","0000001010101101","0000010001001010","0000011010100111","0000100010100101","0000100111000101","0000101100011000","0000110100111101","0000111100011000","0000111101011010","0000111001100111","0000110111100011","0000111011000001","0001000000100111","0001000001010010","0000111010100111","0000110010101101","0000110000101011","0000110001111011","0000101101000010","0000100000001111","0000010101001100","0000010010000111","0000001111010010","0000000011000110","1111110001110011","1111100111011010","1111100110001010","1111100101011101","1111100000001110","1111011001010111","1111010010110100","1111001010111010","1111000011100111","1111000010101100","1111000111010001","1111001000100111","1111000011001110","1110111111000001","1111000011000111","1111001010110111","1111001101101110","1111001100110111","1111010000100110","1111011010101010","1111100011100011","1111100110011100","1111101000111000","1111110010100110","0000000010000011","0000001110011110","0000010100001100","0000011000111111","0000100010100010","0000101101011001","0000110010011000","0000110001110011","0000110011000100","0000111001100011","0000111111111101","0001000000110001","0000111101111100","0000111100101101","0000111101101110","0000111101001111","0000111000101110","0000110001001111","0000101001101101","0000100100011110","0000100001000101","0000011011111000","0000010010011011","0000000111110111","0000000000110111","1111111011101111","1111110010100101","1111100101110010","1111011100110010","1111011001111101","1111010101110111","1111001011011111","1111000001000001","1110111110010010","1111000000110111","1111000001110000","1111000001010000","1111000100010011","1111001001110001","1111001011101011","1111001001010001","1111000111111110","1111001010111110","1111010000100100","1111010111001000","1111011110011010","1111100101100010","1111101100100111","1111110110101001","0000000011111000","0000001110001001","0000010001010001","0000010011011111","0000011100100100","0000101000100011","0000101101101111","0000101101011110","0000110010001110","0000111101000000","0001000010001100","0000111100101101","0000110111000110","0000111011000110","0001000010100101","0001000001101110","0000111000011000","0000110000010001","0000101110001011","0000101101101101","0000101001011000","0000100000010011","0000010100011111","0000001000110100","1111111111101100","1111111000010111","1111101110110101","1111100001110011","1111010110101011","1111010011101100","1111010110111101","1111010111100100","1111010000000001","1111000101000101","1111000000000000","1111000011001000","1111000110011101","1111000001110001","1110111000100110","1110110111011001","1111000011101000","1111010011111001","1111011011110010","1111011011001011","1111011011010110","1111100001000101","1111101001010101","1111110001101000","1111111011010101","0000000110000110","0000001110111011","0000010101111001","0000011110000010","0000100110101000","0000101011101001","0000101101110110","0000110010110101","0000111010111111","0000111111100101","0000111101101000","0000111011000011","0000111100111100","0000111111110101","0000111110000111","0000111000010011","0000110001110101","0000101011001111","0000100100010100","0000011110111011","0000011011000110","0000010100111000","0000001010111010","0000000010001100","1111111110010110","1111111011000111","1111110011000111","1111101000100100","1111100001000100","1111011100001110","1111010101011111","1111001100110100","1111000110100110","1111000100011001","1111000011101110","1111000011011000","1111000100101101","1111000111011110","1111001001100110","1111001010110101","1111001100111000","1111001111101110","1111010001110111","1111010011111100","1111011000101111","1111100001000100","1111101010101011","1111110011001010","1111111010000110","0000000000011010","0000000111111100","0000010010011000","0000011110101100","0000101000110011","0000101110000010","0000110000011010","0000110011011100","0000110111010111","0000111010000000","0000111010110100","0000111011010100","0000111100100011","0000111110011110","0001000000100000","0001000000110011","0000111100101110","0000110100010000","0000101010111001","0000100011011111","0000011100111000","0000010100111011","0000001100001101","0000000100000011","1111111011011100","1111110001001101","1111100111010001","1111100000100011","1111011100111001","1111011001010001","1111010011010101","1111001011000011","1111000010100111","1110111101111000","1110111110111000","1111000010000000","1111000001000110","1110111100010101","1110111011100000","1111000011010111","1111001110011111","1111010100111001","1111010110100100","1111011001011011","1111011111111010","1111100111011111","1111101110101110","1111110111010000","0000000001110110","0000001100101111","0000010101110001","0000011011101101","0000011110101101","0000100001001100","0000100110101101","0000101111011001","0000110111011101","0000111100100110","0001000000100110","0001000100010011","0001000100111100","0001000001110010","0000111110111011","0000111110011100","0000111100000000","0000110100111000","0000101110000100","0000101011101101","0000100111111010","0000011011011010","0000001010111111","0000000010000110","0000000010001001","0000000001100101","1111111010111101","1111110010001001","1111101010000001","1111011111111111","1111010100011111","1111001101100101","1111001100101001","1111001010011001","1111000010011101","1110111010110000","1110111010000011","1110111110000111","1111000001010011","1111000011100100","1111000111000011","1111001001110101","1111001010110100","1111001111101100","1111011101000111","1111101100011000","1111110010100011","1111110000101001","1111110010111000","1111111110100111","0000001010111100","0000001111000011","0000001111101000","0000010110110010","0000100100011000","0000101111000001","0000110010111001","0000110110100011","0000111111011011","0001001000100101","0001001001111110","0001000100011010","0001000000000000","0001000000011100","0001000000110000","0000111011111101","0000110100001000","0000101110000110","0000101001110000","0000100011010100","0000011010001010","0000010001111111","0000001100111010","0000000111110111","1111111110110011","1111110010010111","1111100111100000","1111100001011001","1111011101110011","1111011000001110","1111001111101010","1111000111011001","1111000010001000","1110111111001110","1110111101110101","1110111111011000","1111000100000000","1111000111100111","1111000110111110","1111000101110011","1111001010001010","1111010010110001","1111011000000111","1111011000001011","1111011010010011","1111100100011100","1111110010100110","1111111101010100","0000000011111000","0000001011000111","0000010100110100","0000011101110000","0000100011001101","0000100101111100","0000101000010101","0000101100001001","0000110001111001","0000111000010101","0000111100111001","0000111110001111","0000111101011011","0000111011111001","0000111010000010","0000111000000000","0000110101011001","0000110000000101","0000100110100100","0000011100010010","0000010110110110","0000010101100101","0000010001100110","0000001000000111","1111111110111101","1111111010100100","1111110110001100","1111101011101000","1111011101101100","1111010011111000","1111001111100101","1111001100110101","1111001010001001","1111001000000101","1111000100010101","1110111101101110","1110111010001010","1110111111001111","1111000111010101","1111001000100000","1111000100110100","1111000111110001","1111010011000001","1111011011100001","1111011100110111","1111100001001010","1111101110110111","1111111100010000","1111111111010001","1111111110101111","0000000110110001","0000010100010110","0000011011001000","0000011011000010","0000100000100011","0000101111000101","0000111010011001","0000111001011110","0000110011100010","0000110011110001","0000111001010111","0000111100100001","0000111100000011","0000111100100100","0000111101100010","0000111001011011","0000110000001100","0000101000111011","0000100110110110","0000100100001011","0000011011010111","0000001111001101","0000000100111110","1111111011111000","1111110000110011","1111100110010011","1111100001101001","1111100001011011","1111011110011100","1111010101101100","1111001011001101","1111000010110110","1110111100111110","1110111010100111","1110111110000011","1111000101000101","1111001001001111","1111001000001011","1111000110101001","1111001001000111","1111001110110011","1111010101110001","1111011101111100","1111100101111010","1111101011001110","1111101111110110","1111111000110100","0000000101000010","0000001100101110","0000001101100010","0000001111001010","0000010111011000","0000100001110000","0000101000100010","0000101101110011","0000110100101110","0000111001011000","0000111000010011","0000110111000101","0000111011110101","0001000001001110","0000111110001011","0000110101010010","0000110001000010","0000110010110100","0000110001101000","0000101001100100","0000100000110011","0000011011101000","0000010110010001","0000001101111100","0000000110010011","0000000001100011","1111111011011001","1111110000110111","1111100101111010","1111011110011010","1111010111111101","1111001111101111","1111001000011111","1111000101011001","1111000100010100","1111000010001010","1110111111111100","1110111110111110","1110111101011110","1110111100000001","1111000000001111","1111001011011001","1111010100110000","1111010101010101","1111010100001110","1111011101010001","1111101110111010","1111111011101100","1111111101010000","1111111011111110","0000000001110010","0000001110011010","0000011010111100","0000100010111100","0000100110110101","0000101001110111","0000110000001011","0000111010011101","0001000010111001","0001000010101000","0000111011011100","0000110111000101","0000111011000110","0001000010000010","0001000011010110","0000111101110101","0000110110011111","0000110000010011","0000101001111100","0000100010110011","0000011101000100","0000011001011000","0000010011101001","0000000111101011","1111110111110100","1111101011010011","1111100101100110","1111100010010001","1111011011101000","1111010010001000","1111001010011101","1111000110101111","1111000101011010","1111000101011001","1111000110100010","1111000110110000","1111000011101001","1110111111101111","1111000000111010","1111001000100000","1111010000111111","1111010101100111","1111010111111100","1111011011101000","1111100000100000","1111100100110010","1111101001110101","1111110010010101","1111111100111011","0000000101100111","0000001011111101","0000010011101101","0000011110001101","0000100111011000","0000101011110110","0000101110111010","0000110101110001","0000111110101001","0001000010001001","0000111110100101","0000111011100011","0000111110100010","0001000001111111","0000111101110011","0000110100111011","0000110001011011","0000110100001100","0000110010010000","0000100101000101","0000010100101000","0000001100000010","0000001010101010","0000000111000101","1111111100110011","1111110000000111","1111100110011100","1111100000100111","1111011100001111","1111010110110101","1111001111101101","1111001001001101","1111000110111010","1111001000011101","1111001000111011","1111000101011001","1111000001000101","1111000000000001","1111000001110110","1111000101100010","1111001101001001","1111011000001100","1111011111001010","1111011100110100","1111011000111010","1111011111100101","1111101111011100","1111111011001001","1111111101111011","0000000010010111","0000001111110110","0000011101011111","0000100000110010","0000011111100010","0000100110101011","0000110100110010","0000111100001000","0000111000101110","0000110101101111","0000111010100010","0000111111100101","0000111100110001","0000110111000001","0000110110011000","0000110111101100","0000110011000010","0000101010010100","0000100101100000","0000100011111100","0000011101011011","0000010000110101","0000000110000100","0000000000100111","1111111010110000","1111110000101110","1111100110010111","1111011110101001","1111010110110100","1111001110000111","1111001001110100","1111001100010000","1111001110101101","1111001010011000","1111000001111001","1110111100110001","1110111101111000","1111000011000101","1111001001110011","1111001111101101","1111010010001100","1111010001011111","1111010001101011","1111010110010011","1111011111000101","1111101010001101","1111110101100100","1111111101011111","1111111111010101","1111111111000000","0000000100100001","0000010010001010","0000100001011011","0000101011001111","0000101110110000","0000101111011010","0000110001000101","0000110110101100","0000111111011110","0001000101101010","0001000100111010","0001000001000110","0001000000010101","0001000000011010","0000111010110010","0000110001101000","0000101101110001","0000101110111100","0000101010001100","0000011011011010","0000001100011100","0000000101101010","0000000010000011","1111111001010100","1111101100110110","1111100010101100","1111011011110000","1111010110010100","1111010011101000","1111010011000011","1111001110011010","1111000011100001","1110111011001110","1110111101100111","1111000100100010","1111000100100010","1110111110110100","1110111110111010","1111000111101111","1111010000000101","1111010010100001","1111010101100000","1111011111001011","1111101011001011","1111110010011000","1111110101010000","1111111000110101","1111111111001010","0000000111110111","0000010011011010","0000100000001011","0000101000101100","0000101010100111","0000101011100101","0000110001011010","0000111001000011","0000111011110100","0000111010001111","0000111010100001","0000111110000000","0000111111110101","0000111101110100","0000111011000111","0000111000110001","0000110011000011","0000101001000010","0000100000011010","0000011101010011","0000011010110101","0000010001101001","0000000011100001","1111111001111111","1111111000111110","1111111000101110","1111110000001000","1111100000011110","1111010010101010","1111001011100101","1111001000101011","1111000110110111","1111000110001010","1111000101110001","1111000011010000","1110111111110110","1111000000001010","1111000011111100","1111000101000001","1111000010010001","1111000011110100","1111001110011100","1111011010110010","1111100000111000","1111100100101001","1111101101100101","1111111000110111","1111111111001110","0000000010100111","0000001001110110","0000010011000000","0000010111110101","0000011100000010","0000101000011101","0000111001001100","0001000000001001","0000111010010001","0000110100000110","0000110110011101","0000111100010011","0000111110111011","0000111111101110","0001000000011010","0000111101011110","0000110101111111","0000101111100011","0000101101000000","0000101001100101","0000100001011111","0000010111101001","0000001110101010","0000000100010100","1111111000000010","1111101110000101","1111101000010011","1111100010100111","1111011010101000","1111010100000001","1111010001011011","1111001111100101","1111001011010001","1111000110010010","1111000010111010","1111000000010101","1110111110000011","1110111101101001","1110111111001001","1111000001001011","1111000101100111","1111001111000101","1111011000111101","1111011011000000","1111010111000101","1111011001011100","1111100111001011","1111110110001010","1111111100011110","1111111110110100","0000000111001101","0000010100111100","0000011111011101","0000100100100001","0000101001100111","0000110001011000","0000111000100101","0000111100100000","0000111101110111","0000111101110000","0000111101001101","0000111110011100","0001000001010011","0001000000101001","0000111001100100","0000110010001010","0000110001101110","0000110100001010","0000101110010100","0000011110101110","0000010000011000","0000001010101001","0000000111100011","1111111110100000","1111110000011110","1111100100001001","1111011011111100","1111010110001001","1111010010011010","1111010000111101","1111001111001101","1111001010101111","1111000101011101","1111000010100100","1111000001110010","1111000001100001","1111000010111111","1111000111010000","1111001011001000","1111001011010100","1111001010110111","1111001111111000","1111011010100001","1111100100101111","1111101010111011","1111101111101001","1111110110000001","1111111101001010",
--"0000000011011111","0000001010111010","0000010101111100","0000100010110001","0000101100010000","0000101111111110","0000110001010101","0000110101011000","0000111100011110","0001000001110011","0001000001100101","0000111110010001","0000111101100010","0001000000111000","0001000011100011","0001000000101001","0000111000111011","0000110000111111","0000101011011101","0000100110100101","0000011111000101","0000010011101011","0000000110101010","1111111100011100","1111110111101011","1111110101101100","1111101111110101","1111100010101001","1111010011010100","1111001011010000","1111001101001010","1111010001010000","1111001110011010","1111000101000101","1110111101001011","1110111011000100","1110111011100000","1110111011011000","1110111101000101","1111000011000111","1111001010001101","1111001110011010","1111010010001000","1111011010011001","1111100101111111","1111101110101010","1111110010110000","1111110111010110","1111111111101001","0000001000010011","0000001101100111","0000010010000101","0000011010110100","0000100111011101","0000110001011110","0000110100000001","0000110010010000","0000110011100100","0000111001110011","0000111110100001","0000111100010110","0000110111100110","0000110111111000","0000111011101111","0000111010011110","0000110010100110","0000101100101110","0000101100011011","0000101001000100","0000011011111001","0000001100011011","0000000101001111","0000000011011111","1111111100101000","1111101111100000","1111100100000110","1111011101000100","1111010101100110","1111001101000011","1111001001000001","1111001010000010","1111001000110000","1111000001101001","1110111010110010","1110111010010111","1110111111000010","1111000100111110","1111001011010111","1111010001000100","1111010010110100","1111010001011010","1111010011110110","1111011110011100","1111101011111110","1111110100100001","1111110111100101","1111111011010001","0000000011111101","0000001111111011","0000011001110001","0000011101011110","0000011101010000","0000100000110001","0000101011110001","0000110111000111","0000111001011101","0000110110000100","0000111000111111","0001000011010100","0001000111011010","0000111110000111","0000110011010110","0000110100010110","0000111011100001","0000111010000101","0000101110011101","0000100011011010","0000011101100001","0000010111001011","0000001101110000","0000000101100011","1111111111110110","1111111000011111","1111101110111110","1111100111101100","1111100010010110","1111011001000110","1111001100000111","1111000100000001","1111000100111111","1111000111110110","1111000100110111","1110111110001111","1110111010101001","1110111011011101","1110111101111000","1111000001000010","1111000101101001","1111001011000010","1111010000101000","1111010111011110","1111011111011100","1111100110101001","1111101101100010","1111110111011000","0000000011100101","0000001100001011","0000001110111111","0000010010111100","0000011101111110","0000101010100010","0000101111000010","0000101100111001","0000101110110101","0000111000100101","0001000001101111","0001000011000010","0000111111110001","0000111110000010","0000111101001010","0000111010000111","0000110111000010","0000110110101110","0000110101100111","0000101111010000","0000100111001100","0000100011100100","0000100001010000","0000010111010111","0000000110000011","1111110111110111","1111110010100101","1111101111111111","1111101000111011","1111011110110010","1111010110010011","1111010000011100","1111001100110100","1111001100001110","1111001100010011","1111000111100010","1110111101111001","1110110111011011","1110111001011101","1110111111100001","1111000011100000","1111000110001011","1111001010011111","1111001111000101","1111010010110001","1111011001010111","1111100100111101","1111101111110110","1111110100001101","1111110101110110","1111111100101011","0000001001011010","0000010110100111","0000100001100000","0000101010100101","0000110000001101","0000110000011000","0000101110011101","0000110000010001","0000110110010011","0000111100001110","0000111111110000","0001000001010011","0000111111011011","0000111000110111","0000110001111010","0000110000111001","0000110100000011","0000110001111000","0000100101101010","0000010110011111","0000001110010000","0000001101010011","0000001011000000","0000000000101100","1111110000110100","1111100011000000","1111011011110011","1111011000111011","1111010101000010","1111001101110010","1111000101101001","1111000000011010","1110111111001001","1110111111100100","1110111110111011","1110111101000011","1110111100111010","1111000001000011","1111000111110000","1111001100010001","1111001101001011","1111001110110110","1111010101100001","1111011111010101","1111100111101001","1111101110000100","1111110101010110","1111111101011010","0000000100010010","0000001100010001","0000011001011110","0000101000001110","0000101110100110","0000101010110011","0000101000011000","0000110000101001","0000111100110100","0001000000010000","0000111011011111","0000111010101110","0001000010011101","0001001000111100","0001000101011101","0000111100011000","0000110110100011","0000110011110101","0000101101111000","0000100011011011","0000011000111111","0000010000101001","0000001000100110","0000000001000010","1111111100001101","1111111000100000","1111110001001110","1111100110011111","1111011110001101","1111011010101100","1111010110011101","1111001100110010","1111000001010001","1110111011000100","1110111100000010","1111000000011101","1111000100010101","1111000101100010","1111000011100011","1111000000111111","1111000010101100","1111001010001100","1111010011011100","1111011011001000","1111100011011000","1111101110010101","1111111000001000","1111111011111000","1111111100011101","0000000001100100","0000001100111100","0000011000101001","0000100000001100","0000100101110110","0000101101000110","0000110100110100","0000111001011110","0000111010100100","0000111011010111","0000111110110101","0001000011111000","0001000101111001","0001000010000100","0000111011011111","0000110111110100","0000110111011000","0000110100110001","0000101100111010","0000100011001001","0000011010110111","0000010010101001","0000001000111111","0000000000111001","1111111100010001","1111110110101010","1111101011011111","1111011110010101","1111010110011110","1111010100110100","1111010011111011","1111010000000010","1111001001101010","1111000010101011","1110111101101111","1110111101111011","1111000010000101","1111000011111101","1111000000111101","1110111111000000","1111000011010010","1111001001111101","1111001110010110","1111010100110100","1111100010100111","1111110001101010","1111111000100010","1111111010110110","0000000011111111","0000010011000100","0000011011010001","0000011001010111","0000011001111101","0000100101011110","0000110011011100","0000111000110100","0000110111101011","0000111000001001","0000111011000000","0000111100011011","0000111101010101","0001000000011110","0001000010110110","0000111111111011","0000111001111100","0000110101111000","0000110001110110","0000101000001101","0000011011001010","0000010011101100","0000010011110110","0000010010000101","0000000110011010","1111110101100111","1111101010100000","1111100111110111","1111100110110000","1111100001000010","1111010111011000","1111001101001110","1111000100001011","1110111101110011","1110111100111000","1111000000101000","1111000010100100","1110111101111011","1110110111101011","1110111001010110","1111000011111100","1111001110010110","1111010001110110","1111010010100010","1111011000001100","1111100011001100","1111101101100000","1111110011100001","1111110111011111","1111111101001100","0000000101111000","0000010000001101","0000011001110000","0000100001010010","0000101000001110","0000110000010001","0000110111001010","0000111000100001","0000110101100111","0000110110010000","0000111110000000","0001000101011000","0001000011110110","0000111100100001","0000111001001010","0000111010100111","0000110111100011","0000101011100000","0000011110000011","0000010111100001","0000010101101001","0000010000110101","0000000111010111","1111111101110001","1111110111000111","1111110010001010","1111101100101011","1111100101100010","1111011100100101","1111010011011100","1111001101010000","1111001011001100","1111001010110101","1111001001100100","1111000111011000","1111000101000011","1111000010101001","1111000001111000","1111000101111110","1111001110001001","1111010100011010","1111010101110000","1111010111001001","1111011110001010","1111101000001100","1111101110111000","1111110010000110","1111110111000011","1111111111100010","0000001000111101","0000010010111110","0000011111101010","0000101100100101","0000110011001000","0000110010001110","0000110001001110","0000110101111110","0000111101011101","0001000001111100","0001000011100000","0001000101011010","0001000110011011","0001000010010110","0000111010000101","0000110011111111","0000110010100001","0000110000001000","0000100111110000","0000011101000101","0000010110110111","0000010011111001","0000001100100101","1111111111011011","1111110011110101","1111101101111010","1111100111100001","1111011011010100","1111001111101111","1111001101101011","1111010001001111","1111001110011001","1111000011110111","1110111101001111","1111000000110100","1111000110010100","1111000100101010","1110111111010111","1110111111010100","1111000101110010","1111001101101011","1111010100100101","1111011011000111","1111100000001111","1111100011101000","1111101001011011","1111110100111010","0000000001010111","0000000111101111","0000001001100100","0000001110111101","0000011010001000","0000100100011001","0000101001000000","0000101011101111","0000110001101100","0000111001010110","0000111101101000","0000111101100010","0000111100101010","0000111101110001","0000111111111110","0001000000010101","0000111100101110","0000110101110111","0000101111001000","0000101011001111","0000101000110010","0000100011011100","0000011001010011","0000001100101111","0000000001001101","1111111000010110","1111110010011000","1111101101111100","1111100111010110","1111011011110000","1111001110100010","1111000111010100","1111001000100001","1111001011111111","1111001011011101","1111001000000101","1111000110000100","1111000101010110","1111000011100001","1111000010001000","1111000101000111","1111001100000011","1111010010100111","1111010111010000","1111011100011110","1111100011100010","1111101010100011","1111110000101001","1111110111100000","1111111111100011","0000000110011110","0000001011100010","0000010001100110","0000011010100011","0000100011100000","0000101001001000","0000101101100101","0000110101011100","0000111111010000","0001000011011000","0000111110010001","0000110110110111","0000110101110011","0000111001011100","0000111000110110","0000110001111101","0000101100100111","0000101101011101","0000101101111010","0000100110110110","0000011011110100","0000010100001001","0000001110110011","0000000110010010","1111111100000101","1111110101110110","1111110001011001","1111100111011010","1111011001011110","1111010001100110","1111010010000000","1111010001100010","1111001011001101","1111000101100000","1111000100110111","1111000011011110","1110111101110110","1110111100010111","1111000101101101","1111010000111110","1111010001001110","1111001001001101","1111000110111010","1111001111010000","1111011010011111","1111100011010101","1111101100111110","1111111000101100","0000000001000100","0000000011111000","0000001000000101","0000010100010111","0000100100110010","0000101111100001","0000110000111010","0000101110111011","0000110001110100","0000111011101000","0001000110001011","0001001001001101","0001000011100101","0000111100101001","0000111010101100","0000111010101100","0000110101111100","0000101101010110","0000101000000001","0000100111010001","0000100100000100","0000011010010100","0000001110111010","0000000111001100","0000000001010110","1111111001011110","1111110000001100","1111100111011110","1111011110001110","1111010100010111","1111001110001100","1111001101101100","1111001101001110","1111000111100001","1111000000011010","1110111110010010","1110111111001110","1110111101011110","1110111011000000","1110111110110100","1111000111101111","1111001100111001","1111001100001101","1111001110001011","1111011000010100","1111100101011010","1111101111001001","1111110110110011","1111111111010011","0000000110011001","0000001001111111","0000001110100010","0000011000010111","0000100011100100","0000101001000111","0000101001100011","0000101011011010","0000110001000110","0000110111000001","0000111010101010","0000111101000100","0000111110100011","0000111101101001","0000111010111111","0000111001011101","0000111001000110","0000110110010101","0000101111010101","0000100110101110","0000011111010000","0000011000011010","0000010001000111","0000001010100011","0000000101110100","0000000000110010","1111111000011010","1111101101000111","1111100010010011","1111011010001010","1111010011111011","1111001110011101","1111001010000001","1111000110100111","1111000010101101","1110111101010110","1110111000110101","1110111000110000","1110111101001100","1111000010000011","1111000100101111","1111001000001001","1111010000100001","1111011100011111","1111100101110100","1111101001010100","1111101011001111","1111110010000001","1111111110100011","0000001011011110","0000010011010001","0000010110001000","0000011001011111","0000100010000111","0000101110011011","0000110111100110","0000111001001101","0000110110101001","0000110110110010","0000111011010010","0000111111010111","0000111111000110","0000111100110110","0000111100111110","0000111110111001","0000111101001000","0000110100011111","0000101000110000","0000100000110010","0000011110100001","0000011100111110","0000010110100101","0000001011100101","0000000000000001","1111110101101111","1111101011101011","1111100010001111","1111011011101111","1111011000011001","1111010101101110","1111010010010100","1111001110111011","1111001011010011","1111000110101100","1111000011000111","1111000011011100","1111000101110101","1111000110001001","1111000101100101","1111001001001000","1111001111110000","1111010010101001","1111010001110100","1111010110101101","1111100101100110","1111110101010010","1111111011111110","1111111100100100","1111111111111111","0000000111110001","0000001111110000","0000010111100100","0000100001100100","0000101011110111","0000110010011101","0000110110001011","0000111010110010","0000111111111010","0001000001111111","0001000000110000","0000111111001010","0000111110001111","0000111100111101","0000111011011100","0000111010010000","0000110111011011","0000110000001010","0000100100100011","0000010111100100","0000001100100001","0000000101110111","0000000011011110","0000000000111001","1111111001000001","1111101100101100","1111100001111100","1111011011100100","1111010110100010","1111010000110011","1111001100011101","1111001010000110","1111000110101101","1111000010011100","1111000010010011","1111000110101111","1111001000000110","1111000010011011","1110111110000100","1111000100100100","1111010010001010","1111011011000011","1111011011111111","1111011100101111","1111100011001100","1111101100111100","1111110101110100","1111111101111110","0000000111000100","0000010000110111","0000011001111100","0000100000111110","0000100100110110","0000100111001011","0000101100110100","0000110111011010","0000111111111000","0000111110000101","0000110101011100","0000110010100110","0000111010000101","0001000001011001","0000111101101000","0000110010011110","0000101011110010","0000101100101001","0000101100111010","0000100110101001","0000011101100110","0000010111011010","0000010010110110","0000001010111110","1111111111001011","1111110011101011","1111101011010001","1111100100100010","1111011101001100","1111010101010111","1111001110110110","1111001011000100","1111001001111010","1111001001011111","1111000111010110","1111000011001001","1110111111010101","1110111110000100","1110111110111101","1111000001111100","1111001001010101","1111010100101101","1111011100011010","1111011001110001","1111010011011100","1111011000010111","1111101011100001","1111111110000100","0000000011000100","0000000001000000","0000000110111010","0000010110101100","0000100101000110","0000101011100100","0000101110100011","0000110010011011","0000110100111111","0000110100101000","0000110101011011","0000111011000100","0001000011010100","0001001001100011","0001001011101101","0001001001101010","0001000011010101","0000111001010100","0000101101100100","0000100010110111","0000011100001010","0000011010000110","0000010111111000","0000001110101111","1111111111100110","1111110011110010","1111110000000000","1111101101001111","1111100100110110","1111011011101101","1111011000010010","1111010101000000","1111001001011001","1110111011101110","1110111010001100","1111000011111111","1111001000110111","1111000001101111","1110111010111001","1111000000001101","1111001100010101","1111010011000011","1111010010101100","1111010010100010","1111010110101110","1111011101101110","1111100101111010","1111101110110011","1111110111000001","1111111101101010","0000000100010011","0000001100110111","0000010110111110","0000100000101110","0000101000001101","0000101011111110","0000101101000110","0000110000001110","0000111000001001","0001000000010101","0001000001110000","0000111100111000","0000111000110011","0000111000111001","0000111001101011","0000111000101000","0000110111010100","0000110101011111","0000101111010100","0000100100010111","0000011001110011","0000010010010111","0000001010101000","0000000000011100","1111110111101001","1111110011000101","1111101111001110","1111101000001111","1111100000000010","1111011001110000","1111010100001101","1111001101100010","1111000111111011","1111000101101100","1111000100110000","1111000010011010","1111000000001111","1111000000100001","1111000001111110","1111000011000100","1111000110011000","1111001110010001","1111010111101101","1111011101111010","1111100001010011","1111100110010010","1111101111000101","1111111001111001","0000000011100110","0000001010000001","0000001110000100","0000010100100010","0000100000011100","0000101100000101","0000101110100001","0000101010000100","0000101011110011","0000111000011011","0001000011101010","0001000010011000","0000111011101001","0000111100010100","0001000001111001","0000111111101110","0000110100110100","0000101100110010","0000101011111110","0000101001101011","0000100000011100","0000010110001110","0000010000000010","0000001001111010","0000000000111010","1111111010000010","1111110111111011","1111110011011001","1111100110100011","1111010111101010","1111010000001001","1111001110100000","1111001010100100","1111000010101011","1110111100001111","1110111001111010","1110111010001001","1110111101000001","1111000011001010","1111001000101010","1111001001010010","1111001000111000","1111001111001111","1111011011111010","1111100101110100","1111101000110100","1111101011010100","1111110011110011","1111111111110011","0000001001000010","0000001110101110","0000010100111010","0000011101110010","0000100111110110","0000110000011011","0000110101100110","0000110111000100","0000110111010100","0000111010001111","0001000000100110","0001000110001100","0001000110001001","0001000000101011","0000111011001001","0000111010100101","0000111110000101","0000111110100111","0000110101101111","0000100101100011","0000010111011011","0000010001100001","0000001111110010","0000001010100010","0000000000110110","1111110111101010","1111110000110010","1111101001000100","1111011111100110","1111011000001011","1111010100100000","1111010000101110","1111001001100001","1111000001111001","1110111111000100","1111000001001101","1111000011101011","1111000011000010","1111000000001110","1110111110101110","1111000001001010","1111000111100000","1111001111010110","1111010110111111","1111011111110011","1111101011100101","1111110111111011","1111111111100010","0000000001100100","0000000011111111","0000001100001101","0000010111110011","0000100000010011","0000100100001101","0000101000001010","0000101111001010","0000110101111101","0000111000001110","0000110111100110","0000111010000011","0001000001011110","0001000111111111","0001000110110001","0000111110111101","0000111000100010","0000110111111100","0000111000001000","0000110001111001","0000100110001101","0000011100011001","0000010111010010","0000010010000010","0000001000110010","1111111110000011","1111110100011111","1111101001110000","1111011100101011","1111010011000110","1111010001111010","1111010011011000","1111001101111101","1111000011010100","1110111110110010","1111000100001111","1111001010010000","1111001000010011","1111000001111000","1110111110101000","1110111111010111","1111000001000011","1111000100111110","1111001110001100","1111011010011000","1111100011111101","1111101001110000","1111101111001101","1111110110010111","1111111110010001","0000000101111100","0000001100111111","0000010010100011","0000010111001011","0000011101111111","0000101000100001","0000110011010101","0000111010000010","0000111100101101","0000111110011110","0001000000101011","0001000010011010","0001000010111000","0001000001011101","0000111101110000","0000111001011001","0000110110111000","0000110100101001","0000101101110101","0000100010010000","0000011000010010","0000010011010110","0000001110101110","0000000110001101","1111111101100100","1111111001000110","1111110100111001","1111101011011100","1111100000000010","1111011001101010","1111010111001011","1111010010000111","1111001010010111","1111000101010000","1111000010111000","1110111110100100","1110111001100001","1110111010100100","1111000010010011","1111001001010111","1111001100011001","1111001111111001","1111010110000001","1111011010001000","1111011010101010","1111011101111010","1111100111101101","1111110010100001","1111111001011000","0000000000100101","0000001100111011","0000011001001101","0000011110000101","0000011111000001","0000100101000001","0000101111100100","0000110110010000","0000110111110000","0000111011100000","0001000011010001","0001000110111010","0001000010011111","0000111101101111","0000111111000111","0001000000111000","0000111010110111","0000101111101011","0000100111010100","0000100010101011","0000011101011001","0000010111011101","0000010010110011","0000001011100111","1111111101101011","1111101110011110","1111100110101101","1111100011101011","1111011011100000","1111001110100101","1111000111011101","1111001000010101","1111000111011100","1111000001010001","1110111111010100","1111000110011000","1111001100001001","1111001000001100","1111000010011011","1111000101101011","1111001110001110","1111010010010110","1111010011100011","1111011001010110","1111100001101001","1111100101001001","1111100111010111","1111110010011011","0000000100011100","0000010000000000","0000010001001001","0000010011101111","0000100000101001","0000110000011111","0000110111111101","0000110111110100","0000111001000001","0000111110111000","0001000100101100","0001000110000000","0001000010110111","0000111101110001","0000111001100011","0000111000100000","0000111001111110","0000111001010101","0000110010100101","0000100111100101","0000011110001001","0000011000100111","0000010011001100","0000001010010001","0000000000011001","1111111010010101","1111110110010000","1111101100111100","1111011101101101","1111010010100110","1111010010110011","1111010110010100","1111010000001111","1111000010011000","1110111011011110","1111000001110000","1111001011000010","1111001100110100","1111001001010100","1111000111010110","1111000111110101","1111001010010110","1111010010000000","1111011110010000","1111100111000001","1111101000001110","1111101001010011","1111110000110110","1111111010001000","1111111111101100","0000000111000010","0000010101110000","0000100011110101","0000100110110111","0000100100010000","0000101001010111","0000110110001101","0000111111011000","0001000001101110","0001000100000001","0001000110111100","0001000011101001","0000111011010000","0000110111011110","0000111001010111","0000110110101111","0000101100001100","0000100011010101","0000100010000001","0000100000110111","0000011000011101","0000001100010111","0000000010011011","1111111001110111","1111110001100101","1111101101000101","1111101011110101","1111100101101011","1111010111100110","1111001011011010","1111001010000001","1111001101011110","1111001010011101","1111000001101011","1110111101010000","1111000000001110","1111000011100111","1111000011000011","1111000010111010","1111000111101000","1111001110101100","1111010011100100","1111010110110001","1111011100001111","1111100101011010","1111101111110100","1111111000100111","1111111111011100","0000000101111101","0000001101010110","0000010101000101","0000011100000111","0000100010101011","0000101001101000","0000110000001111","0000110100010101","0000110101111000","0000111000100101","0000111111000001","0001000101110001","0001000110101101","0001000001000111","0000111010110110","0000111000010000","0000110111000010","0000110010111111","0000101100001000","0000100100011110","0000011011100010","0000010000110110","0000001000001100","0000000100110100","0000000010011101","1111111001111100","1111101100011101","1111100010010111","1111011110000100","1111011000111100","1111001111111101","1111001001100100","1111001001110000","1111001001010101","1111000001011111","1110111000110011","1110111010000001","1111000010111101","1111000111110111","1111000101100101","1111000100111100","1111001011010110","1111010011011011","1111010111110001","1111011011100011","1111100011010011","1111101101010001","1111110101111100","1111111110010011","0000001000001101","0000010001011000","0000010111010010","0000011011110010","0000100001010010","0000100110001110","0000101001011000","0000101110111001","0000111010011001","0001000110111100","0001001011101111","0001000111111111","0001000011011001","0001000010010100","0001000000011011","0000111001010111","0000110000110000","0000101100110001","0000101100011010","0000101001000100","0000100000010100","0000010110011110","0000001110010000","0000000100010001","1111110110010111","1111101010100100","1111100111101110","1111101010000101","1111100110111111","1111011100000110","1111010010010011","1111001111000100","1111001100100001","1111000100111111","1110111101100011","1110111100011110","1110111101100101","1110111010001100","1110110110111010","1110111100101100","1111001000100100","1111001111011100","1111010000111001","1111010111011101","1111100101100001","1111110000010011","1111110001111011","1111110011000010","1111111100001011","0000001001001010","0000010010011101","0000011000110111","0000100000001011","0000100110100110","0000101001111101","0000101110010011","0000110111000010","0000111111010010","0001000001000011","0000111110111010","0000111111000100","0001000000110110","0000111111010110","0000111010101101","0000110111001101","0000110101001110","0000110000110100","0000101000101001","0000011111010110","0000010111001000","0000010000010100","0000001011001000","0000000110100101","1111111111010110","1111110011111111","1111101000110000","1111100010100001","1111011111000111","1111010111110000","1111001011001100","1111000000010001","1110111100111010","1110111110110001","1110111111110001","1110111110101100","1110111111000010","1111000001101110","1111000011001110","1111000010011100","1111000100011101","1111001101100000","1111011001111101","1111100011000100","1111101000001000","1111101101000111","1111110010101001","1111110110110001","1111111100001001","0000000111010000","0000010100010010","0000011010011110","0000011010111000","0000100000100011","0000101110010011","0000111000110001","0000111000100010","0000110110000100","0000111010110110","0001000010001000","0001000011001010","0001000000100001","0001000001001001","0001000010011001","0000111101111011","0000110110010100","0000110001011010","0000101100001100","0000100001010001","0000010101100010","0000010000100110","0000001110000010","0000000100100011","1111110111011010","1111110001000001","1111101111100110","1111100111110001","1111011001100000","1111010001000111","1111010010001000","1111010001110101","1111001010010100","1111000011110001","1111000100110010","1111000111100001","1111000100111100","1111000000000111","1110111110110001","1111000000001010","1111000010000101","1111000110111010","1111010000001110","1111011010010001","1111100001111100","1111101001100010","1111110010111000","1111111010111011","0000000000010001","0000000111010101","0000010010111110","0000011110011011","0000100100100011","0000101000001000","0000101110011001","0000110101101101","0000111000011110","0000110110111010","0000110111000100","0000111011011000","0000111111011110","0000111111100001","0000111101011101","0000111100101111","0000111100001111","0000110111110100","0000101110110100","0000100101111010","0000100001100001","0000100000001111","0000011100110110","0000010100101011","0000001001101101","1111111110010111","1111110010101000","1111100110110010","1111011101101010","1111011001000100","1111010101111011","1111001111111011","1111000111111111","1111000011000111","1111000011000011","1111000011111110","1111000010011111","1110111111111001","1110111110111101","1111000000000110","1111000010111110","1111001000101101","1111010001001010","1111011000110000","1111011100111101","1111100001010010","1111101011000110","1111111001000111","0000000100000010","0000001000101001","0000001100001001","0000010100010001","0000011111000100","0000100110100001","0000101001011100","0000101100011101","0000110010111010","0000111010101000","0000111111010100","0000111111010010","0000111100010100","0000111001011000","0000111000010010","0000111000110111","0000111001100011","0000111000110000","0000110101000101","0000101101011010","0000100010110011","0000011001101010","0000010101100001","0000010011100100","0000001101100011","0000000010111000","1111111001100001","1111110011110111","1111101100001100","1111011110111010","1111010010010001","1111001101000010","1111001011100010","1111000110011101","1111000000000011","1110111111101011","1111000011100011","1111000010111111","1110111101111011","1110111101101101","1111000100111100","1111001011010010","1111001100110100","1111010000100011","1111011010000101","1111100001110111","1111100011100010","1111100111011000","1111110011100001","1111111111011000","0000000010001110","0000000100000110","0000010001000111","0000100011100000","0000101011011001","0000101000001000","0000101000100000","0000110010010011","0000111011010011","0000111100100111","0000111100101110","0001000000111011","0001000011100011","0000111111110100","0000111011010111","0000111011001110","0000111010000111","0000110010000011","0000100111000110","0000011111111000","0000011010111100","0000010100010010","0000001110000000","0000001010011001","0000000100000110","1111110110010011","1111100111010111","1111100000111001","1111100001001110","1111011110110101","1111010110110011","1111001101111000","1111000110010000","1110111110110100","1110111010100000","1110111101001000","1111000010000111","1111000001110011","1110111111000111","1111000011101101","1111001110110001","1111010101010000","1111010100101110","1111010111101111","1111100010101111","1111101011111110","1111101101001100","1111101111011100","1111111010111101","0000001000000100","0000001100100100","0000001101110010","0000010110110001","0000100100010111","0000101010110000","0000101010010100","0000101111000001","0000111100001000","0001000110111100","0001000111011111","0001000001111110","0000111101010011","0000111010001110","0000110111011111","0000110101110111","0000110100110100","0000110001101101","0000101100010010","0000100110100100","0000011111111010","0000010110010011","0000001100001010","0000000101100000","1111111111101001","1111110100001101","1111100100110100","1111011010101101","1111011000100110","1111010110011111","1111001110110011","1111000111011000","1111000111100000","1111001011111101","1111001011111110","1111000110001011","1111000001101001","1111000011011010","1111001000011101","1111001011001010","1111001011000011","1111001100110111","1111010011100010","1111011011101101","1111100000110001","1111100100011001","1111101100100101","1111111010000001","0000000110001100","0000001101001100","0000010010111111","0000011010101111","0000100000010011","0000100000110010","0000100010111010","0000101101011001","0000111010001001","0000111101110101","0000111001100011","0000111000110111","0000111111000010","0001000010101001","0000111110001110","0000111001010011","0000111010111001","0000111101010101","0000110111010010","0000101010010011","0000011111111000","0000011011110000","0000011000110111","0000010010000100","0000000111111111","1111111101110110","1111110101010110","1111101110001101","1111100111100000","1111100000100110","1111011001101101","1111010011010000","1111001100110011","1111000110001110","1111000001100111","1111000001001101","1111000010111001","1111000001101111","1110111101100001","1110111100011110","1111000010110110","1111001100011101","1111010010100011","1111010101000010","1111011001001011","1111100000111011","1111101001001000","1111110000001001","1111111000111001","0000000101100000","0000010010110000","0000011011101100","0000011111101110","0000100010101111","0000101000001001","0000101111011111","0000110101011001","0000110111011000","0000110110101110","0000110111011011","0000111011010001","0000111110101100","0000111101000110","0000110111110101","0000110100110110","0000110101110110","0000110101011010","0000101111110101","0000101001011111","0000100111010010","0000100100101001","0000011001011001","0000001000000111","1111111100110100","1111111011101010","1111111010010011","1111101111100100","1111100001010101","1111011010100011","1111011001100111","1111010011100100","1111000110010110","1110111100010000","1110111100000101","1110111111111111","1111000000001100","1110111110110010","1111000010011100","1111001010100011","1111001111100100","1111001101101101","1111001001110100","1111001011011000","1111010100011001","1111100000001100","1111101001010001","1111101111100101","1111110111101010","0000000011000001","0000001100110000","0000010000111110","0000010100010111","0000011101110100","0000101010011110","0000110000101110","0000101111011100","0000110000110100","0000111010100001","0001000100001100","0001000100011011","0000111110101111","0000111100001000","0000111100010001","0000111000100110","0000110001110100","0000101110111110","0000101111110000","0000101011110111","0000100001001100","0000010111110011","0000010011111000","0000001110001010","0000000000110100","1111110010100111","1111101100101001","1111101011101000","1111100110000000","1111011100001001","1111010110100011","1111010101110110","1111010001000100","1111000101111011","1110111110101100","1111000010011010","1111001001101101","1111001010101101","1111000111110011","1111001001010100","1111001111000001","1111010010001110","1111010010011111","1111010101100001","1111011100011100","1111100011000111","1111101001000100","1111110001100011","1111111010111100","0000000000100010","0000000100111110","0000010000010101","0000100001101001","0000101101101101","0000101111110011","0000110000011110","0000110110010101","0000111011001100","0000111000011111","0000110100010001","0000110111011000","0000111101110100","0000111101000010","0000110101101001","0000110010010010","0000110110001010","0000111000001000","0000110001001110","0000100101110110","0000011101000001","0000010110100001","0000001110111010","0000000111001011","0000000001111101","1111111101001100","1111110100101010","1111101001100100","1111100001100101","1111011101111110","1111011001010111","1111010000001101","1111000110111101","1111000011100011","1111000100001111","1111000010001101","1110111100101101","1110111011001101","1111000010100100","1111001101010111","1111010011000000","1111010010110010","1111010011010011","1111011000011101","1111011111011001","1111100100011101","1111101000101111","1111101111111110","1111111011010011","0000000111111111","0000010010110010","0000011011000110","0000100010100000","0000101001010011","0000101101010000","0000101101011001","0000101101100101","0000110010111100","0000111100110100","0001000100101010","0001000101111111","0001000010100101","0000111101110011","0000111000110110","0000110101001011","0000110101000110","0000110110100000","0000110010011001","0000100110100111","0000011010101001","0000010101000111","0000010001101001","0000001000100111","1111111100010111","1111110101000011","1111110001111111","1111101010000111","1111011011011110","1111001111100111","1111001101000111","1111001110011011","1111001011110000","1111000110001111","1111000011010000","1111000010110100","1111000001010110","1110111111001110","1111000000011111","1111000110011101","1111001110000110","1111010011110110","1111010110010101","1111010110111110","1111011001100001","1111100000111101","1111101011100001","1111110100011011","1111111010011100","0000000001001010","0000001010110110","0000010101000001","0000011100111100","0000100011000000","0000100111111110","0000101011010001","0000101110001000","0000110011100011","0000111011000011","0000111111110100","0000111111101011","0000111110001111","0000111110000101","0000111100001000","0000110101100100","0000101101101111","0000101001011100","0000100111111101","0000100101001001","0000011111010101","0000010111001110","0000001100110100","0000000000101111","1111110110011110","1111110000110100","1111101101010001","1111100110110110","1111011100110111","1111010011100010","1111001110100000","1111001101000110","1111001100001101","1111001001110110","1111000101111110","1111000001010010","1110111100111000","1110111011000100","1110111110101000","1111000111001010","1111001111001000","1111010001010101","1111010000001100","1111010011100000","1111011101111000","1111101001101011","1111110010000000","1111111000101100","0000000000000010","0000000101101001","0000001000111111","0000010000000110","0000011110010010","0000101100000100","0000110001010011","0000110010001000","0000110111111101","0001000001011100","0001000100111011","0001000000111100","0000111110001010","0001000000011110","0001000001101001","0000111101011011","0000111000000111","0000110101000111","0000110000011011","0000100111000010","0000011101101010","0000011000111011","0000010100111011","0000001011010100","1111111101101101","1111110011010111","1111101110111011","1111101100001011","1111100111001100","1111100000011011","1111011001010000","1111010001001010","1111001000100110","1111000011010000","1111000011111101","1111000111100000","1111000111011001","1111000010010000","1110111110000001","1110111111110100","1111000101011000","1111001001101100","1111001100111011","1111010010100110","1111011010001101","1111100000000001","1111100100011010","1111101011111001","1111110111000110","0000000001001100","0000000111010110","0000001100010111","0000010011011101","0000011100101111","0000100111100110","0000110010101100","0000111001001110","0000110111101100","0000110100000100","0000111000100000","0001000011100110","0001001000000101","0001000000100101","0000111000101100","0000111011001101","0001000001000111","0000111100110010","0000101110100100","0000100010000101","0000011011110000","0000010101010101","0000001011010110","0000000010000101","1111111100100110","1111111000001001","1111110010001110","1111101011101100","1111100100101010","1111011100001000","1111010100001001","1111001111101100","1111001100101110","1111000111000110","1111000000110101","1110111111001001","1111000000010011","1110111101111000","1110111001101101","1110111101000101","1111001000101000","1111010000110001","1111001111010100","1111001101011001","1111010100100011","1111100000010001","1111100111101011","1111101100111000","1111110111101111","0000000111000110","0000010010101011","0000011000010001","0000011101000010","0000100011100000","0000101001011011","0000101110000100","0000110010100001","0000110101010100","0000110100110000","0000110100001010","0000110111100001","0000111011111110","0000111100010101","0000111010001101","0000111010101000","0000111011110010","0000110111101010","0000101111011001","0000101010000100","0000101000000111","0000100010000100","0000010101000010","0000000111001001","1111111101110100","1111110111110011","1111110010110010","1111101110011110","1111101000010001","1111011100111011","1111010000110001","1111001101001000","1111010010010010","1111010101000011","1111001110001101","1111000011111000","1110111110100001","1110111110001000","1111000000000000","1111000110001010","1111010000100010","1111010111000110","1111010100101000","1111010001011001","1111011000100011","1111100111000010","1111110000001101","1111110001001110","1111110011111110","1111111110110111","0000001100011001","0000010101010111","0000011010000101","0000011110101001","0000100100111001","0000101101010001","0000110111001101","0000111110111101","0001000000110011","0000111111100101","0001000001011010","0001000101001000","0001000011011000","0000111011011101","0000110110010100","0000111000111001","0000111100011110","0000111000111011","0000101111000001","0000100011010110","0000010111001110","0000001011101000","0000000100000001","1111111111111010","1111111001000011","1111101101111100","1111100110001001","1111100101011001","1111100011000101","1111010111010000","1111001000100100","1111000010011110","1111000011110101","1111000010101011","1110111101011010","1110111100001000","1111000010001000","1111001001011110","1111001101011001","1111001111110000","1111010011000011","1111010110011111","1111011001011101","1111011101010011","1111100010111010","1111101010011101","1111110100011000","1111111110101000","0000000100001111","0000000100101001","0000000111110100","0000010100101011","0000100110011111","0000110010100010","0000110101100010","0000110100111000","0000110101000101","0000110110011111","0000111001011011","0000111110000110","0001000001110010","0001000010000011","0001000001000011","0001000000111110","0000111110011000","0000110110000001","0000101100001101","0000100110010110","0000100000111110","0000010101111101","0000001001001111","0000000011111100","0000000100001000","1111111101111101","1111101110010110","1111100000000111","1111011010111110","1111011000110111","1111010010000100","1111001001111111","1111001000001110","1111001011001110","1111001010110000","1111000100000111","1110111100101110","1110111010001000","1110111100100001","1111000000111101","1111000101000010","1111001000110101","1111001110100100","1111010111101100","1111100001100111","1111100111110101","1111101010011101","1111101111001100","1111111001101011","0000000110010011","0000001111110011","0000010110101100","0000011110110001","0000100111110010","0000101101111100","0000110000111010","0000110100111110","0000111100001100","0001000010111100","0001000101000111","0001000011010011","0001000000100000","0000111101110011","0000111010101010","0000110111101001","0000110101001010","0000110001010000","0000101001011011","0000011110100111","0000010100101011","0000001110010001","0000001010101100","0000000110101100","1111111110011101","1111110000101100","1111100010000011","1111011010100110","1111011100001110","1111011110010110","1111010111111010","1111001011001110","1111000001111110","1110111110111111","1110111100000010","1110110110000111","1110110011001001","1110110111111100","1111000000011011","1111000110100100","1111001011001101","1111010001110110","1111011001001111","1111011110000111","1111100001111100","1111101000111100","1111110011101100","1111111111010010","0000001001011101","0000010000110111","0000010100101000","0000010111101110","0000011111110101","0000101100010111","0000110011111000","0000110001010100","0000101101110000","0000110100000001","0000111111101101","0001000011101000","0000111110001100","0000111010010001","0000111100010011","0000111100001100","0000110100111110","0000101101011111","0000101011110011","0000101011000110","0000100101000011","0000011100000111","0000010101011011","0000010000001100","0000001001111110","0000000100000110","1111111110010101","1111110011101000","1111100011100111","1111010111011100","1111010101000101","1111010101001111","1111001111011101","1111001000100010","1111001001000010","1111001100101101","1111001000110001","1110111110110110","1110111010101011","1110111110111100","1111000011001110","1111000101001011","1111001100011111","1111011010101000","1111100100111001","1111100100110011","1111100010111000","1111101001100000","1111110101111010","1111111110101101","0000000010110100","0000001001011010","0000010110000000","0000100100000011","0000101101100010","0000110001001001","0000110010000111","0000110100010110","0000111000111010","0000111101001101","0000111110100000","0000111101010011","0000111011111101","0000111011001101","0000111010110000","0000111010111000","0000111010010101","0000110100110110","0000101000110010","0000011100010001","0000010110100000","0000010101001101","0000001111100100","0000000011011111","1111110111111111","1111110001010100","1111101010111010","1111100000101110","1111010110110111","1111010010010100","1111010000010010","1111001011011101","1111000101010110","1111000011000011","1111000011100000","1111000001001001","1110111100001001","1110111011010011","1111000001010010","1111001000101000","1111001100110100","1111010000110010","1111011000000101","1111011111110101","1111100100000010","1111100111101000","1111110000000101","1111111011101101","0000000011111010","0000000111111000","0000001101110001","0000011000000001","0000100001011010","0000100110001010","0000101010100000","0000110011011010","0000111101110111","0001000010110101","0001000001100111","0001000000001001","0001000001101110","0001000010101010","0000111110111000","0000111000110011","0000110110000010","0000110110110011","0000110100101111","0000101011101110","0000100000011001","0000011010001000","0000011000010101","0000010011011000","0000000111110010","1111111010110000","1111110001001011","1111101000100010","1111011101011110","1111010011100111","1111010000001010","1111010000001001","1111001011111011","1111000010101001","1110111011000101","1110111001001101","1110111010000100","1110111011000001","1110111110000000","1111000100000011","1111001001011110","1111001011010111","1111001101001010","1111010100011000","1111100001000101","1111101101110101","1111110110000011","1111111010001110","1111111101101000","0000000010100010","0000001001010000","0000010001110101","0000011100010001","0000100110110110","0000101110000100","0000110000100011","0000110001100101","0000110101001101","0000111010011110","0000111100111000","0000111011000111","0000111000110001","0000111000100001","0000111001000000","0000111000011001","0000110111000100","0000110100101110","0000101111010001","0000100110111111","0000011111101000","0000011010101010","0000010100000000","0000001000011011","1111111011110100","1111110100101001","1111110010111110","1111110000001111","1111100111011100","1111011001111101","1111001100111110","1111000100110111","1111000010101100","1111000011111101","1111000100010101","1111000001101011","1110111110000011","1110111100111000","1110111110110100","1111000010000000","1111000101011011","1111001001101011","1111001110101010","1111010011001010","1111010111101110","1111011111100010","1111101100001110","1111111010000011","0000000011001110","0000000111001001","0000001011010101","0000010011111000","0000011110001101","0000100101100000","0000101001101010","0000101101110100","0000110010010010","0000110101000011","0000110110110101","0000111010100100","0000111111011100","0001000001011001","0001000000000000","0000111111000000","0000111110011011","0000111000110111","0000101100100110","0000100000100100","0000011011100010","0000011010100110","0000010101101001","0000001010011001","1111111101111111","1111110101100111","1111110001010100","1111101101011111","1111100110111101","1111011101100000","1111010011111100","1111001100110010","1111000111100011","1111000011001001","1111000001000011","1111000010011101","1111000011110001","1111000000100100","1110111011100000","1110111011101010","1111000001111100","1111001000001000","1111001011011001","1111001111111001","1111010111111010","1111011111100101","1111100100110001","1111101011100001","1111110110000111","0000000000001000","0000000110011011","0000001100111101","0000010111000111","0000100000110110","0000100110001000","0000101010111110","0000110100010001","0000111101111110","0001000000100010","0000111101000010","0000111011011110","0000111110110011","0001000010011000","0001000010101000","0001000001000111","0000111111100011","0000111100011111","0000110110100001","0000101110111001","0000100111010010","0000011111101100","0000010111011111","0000001110100000","0000000101000110","1111111011111000","1111110011001010","1111101010010111","1111100001010000","1111011001100100","1111010100111000","1111010001001111","1111001011101000","1111000101100101","1111000011010111","1111000100010100","1111000011010000","1111000000000100","1111000001011001","1111001001011010","1111010000100001","1111010000101011","1111001110101010","1111010001011110","1111010111001110","1111011011010000","1111100001000111","1111101110100110","1111111110110101","0000000110111011","0000000110100111","0000001000111010","0000010011010101","0000011111000101","0000100101011001","0000101000110100","0000101110010010","0000110100110111","0000111001110011","0000111101100000","0000111111111100","0000111101111000","0000110111010001","0000110011001110","0000110111000101","0000111101010000","0000111011011001","0000101111111110","0000100011111011","0000011110110000","0000011110001110","0000011010111010","0000010001101110","0000000110000101","1111111100011101","1111110101001010","1111101101110101","1111100110000111","1111100000000001","1111011011111100","1111010111100000","1111010001101000","1111001100001110","1111001000001011","1111000011010000","1110111101001010","1110111010001000","1110111101000110","1111000010101100","1111000110100101","1111001001110110","1111001111001101","1111010101000100","1111011001001001","1111011101111111","1111100110010101","1111101110110100","1111110100001110","1111111011011101","0000001010001000","0000011010100101","0000100010001001","0000100001100110","0000100011110110","0000101100110111","0000110101011101","0000111001001001","0000111011111101","0001000000000110","0001000001010010","0000111110011111","0000111101100101","0001000000010101","0000111111110100","0000111000001110","0000101111110100","0000101100010100","0000101010000010","0000100011110000","0000011011011001","0000010100010111","0000001100111101","0000000011011100","1111111010110001","1111110100001000","1111101011011100","1111100000011000","1111011001111110","1111011010001110","1111010111111111","1111001101110101","1111000100111010","1111000101111110","1111001000111010","1111000001111011","1110110111100010","1110111001111100","1111001000010011","1111010001001001","1111001110000000","1111001011110011","1111010011111110","1111011110011000","1111100010001100","1111100101011001","1111110000010101","1111111101101001","0000000011111101","0000000111000000","0000010001010001","0000100000111100","0000101001110001","0000101000100110","0000101000000101","0000101111101100","0000111001110000","0000111110011100","0000111111001111","0001000001001101","0001000011001011","0001000001000111","0000111100111111","0000111100011100","0000111111000110","0000111101101110","0000110011110010","0000100101011110","0000011010010110","0000010101001011","0000010010100000","0000001101011011","0000000100001100","1111111001001001","1111101111110011","1111101001010100","1111100011110000","1111011100111110","1111010101011110","1111001111100001","1111001011111110","1111001001010010","1111000101010000","1110111111101001","1110111011001010","1110111011000101","1110111111010010","1111000011110111","1111000110010001","1111001001000011","1111001111010001","1111010110101010","1111011011001111","1111011111011101","1111101001100101","1111111000101010","0000000011110111","0000000111010110","0000001010000010","0000010010101001","0000011101111101","0000100101100111","0000101001101110","0000101101101110","0000110001110101","0000110101111110","0000111101000110","0001000110001100","0001001000001111","0000111110101001","0000110100001001","0000110110010010","0001000001010000","0001000100011001","0000111001111011","0000101101001000","0000100111011111","0000100011110011","0000011001100000","0000001011010110","0000000010100000","0000000000011000","1111111101000000","1111110010100100","1111100100111010","1111011011111101","1111011001011111","1111010111001100","1111001111100101","1111000110000001","1111000001110100","1111000010111001","1111000001110011","1110111100010011","1110111010000101","1111000000010110","1111001000011011","1111001010000110","1111001001011001","1111010000001000","1111011101001011","1111100101010101","1111100100100011","1111100011111110","1111101100010010","1111111010110011","0000000111100100","0000010000001111","0000010111100110","0000011111000110","0000100101011011","0000101010000110","0000101110011100","0000110011110101","0000111010010110","0001000000011001","0001000011010101","0001000001011100","0000111100001110","0000110110110111","0000110010101101","0000101110111011","0000101011101010","0000101010100101","0000101011010110","0000101001111101","0000100011010001","0000011001010011","0000010000101001","0000001010000000","0000000001101110","1111110110000101","1111101010110010","1111100011110101","1111011111010011","1111011000011000","1111001111000111","1111001000101110","1111000111110000","1111001000011001","1111000110011010","1111000010100110","1111000000001000","1111000000000110","1111000010011101","1111000111101001","1111001110010100","1111010010101010","1111010011100111","1111010101010000","1111011010100101","1111100000111110","1111100110000010","1111101101000101","1111111000111101","0000000101001100","0000001100011001","0000010001101010","0000011011001101","0000100110101100","0000101100101000","0000101101110111","0000110010101011","0000111100000111","0001000001100101","0000111111101111","0000111110011110","0001000010111111","0001000110010010","0001000001001011","0000111000100001","0000110100011110","0000110010101010","0000101011000010","0000011101111111","0000010011000011","0000001100010100","0000000101100011","1111111110101111","1111111100100000","1111111101001001","1111110111100010","1111101000100111","1111011000111111","1111010000101011","1111001100110100","1111000111100000","1111000010101011","1111000011101101","1111001000101110","1111001010101111","1111001000000100","1111000101010101","1111000100111000","1111000100101010","1111000100110100","1111001001011101","1111010100001111","1111100000101001","1111101000111111","1111101011110001","1111101011110100","1111101101101110","1111110101101111","0000000100011010","0000010100100011","0000011111011100","0000100011101110","0000100101111100","0000101010011011","0000110001001101","0000110111110100","0000111100000010","0000111100110110","0000111011001110","0000111010000010","0000111010111011","0000111011110110","0000111001111111","0000110101101101","0000110001010101","0000101101010110","0000101000100010","0000100010101000","0000011011111001","0000010011011001","0000001000111100","1111111111000101","1111111000001110","1111110010111110","1111101100110011","1111100110011010","1111100001010101","1111011011010001","1111010001001000","1111000110000010","1111000001001101","1111000011101000","1111000101111010","1111000010101010","1110111101101110","1110111101011001","1111000000111100","1111000011001110","1111000100001011","1111001000110000","1111010001110111","1111011001111100","1111011101101000","1111100001010100","1111101010010100","1111110111010011","0000000011110101","0000001111000110","0000011001101101","0000100000101000","0000100001001111","0000100000010011","0000100101010010","0000101111010100","0000110110011110","0000111000001010","0000111001111011","0000111110110000","0001000010000110","0001000000010110","0000111100110101","0000111011010000","0000111001101001","0000110100111010","0000101110010111","0000101000101001","0000100011000111","0000011011110000","0000010010010001","0000000111101001","1111111101101101","1111110111010110","1111110100101101","1111101111110010","1111100010111010","1111010010110111","1111001010101000","1111001100001110","1111001101111001","1111001000110010","1111000001110000","1110111111101010","1111000000101001","1110111110111110","1110111011000001","1110111010001001","1110111110101100","1111000101111001","1111001100010101","1111010001001010","1111010110011110","1111011111001100","1111101011100100","1111110111101001","1111111111101011","0000000100111011","0000001011011110","0000010100011110","0000011101111100","0000100110011111","0000101101111010","0000110011100000","0000110111111000","0000111101001101","0001000010011011","0001000010001011","0000111011011101","0000110110001100","0000111000001110","0000111011010111","0000110110110100","0000101101011111","0000101000110000","0000101000111011","0000100110100001","0000100000011100","0000011011110111","0000010111100100","0000001100111011","1111111110001100","1111110101100110","1111110011101011","1111101101010011","1111011111001010","1111010100010110","1111010011001100","1111010010000011","1111001000110111","1111000000000110","1111000001111000","1111000111101100","1111000101001111","1110111101010101","1110111100100001","1111000100000101","1111001001111101","1111001011000110","1111001111001010","1111011001010011","1111100011000110","1111101000110000","1111101110101100","1111110111101111","1111111111110011","0000000100001111","0000001000111011","0000010001000011","0000011010001000","0000100001100100","0000101000100101","0000101111101011","0000110100011011","0000110110100101","0000111001100110","0000111110100001","0001000001110010","0001000001001101","0000111110101011","0000111011010011","0000110101110000","0000101111010111","0000101100001110","0000101011111110","0000101000111101","0000100000111101","0000011000100101","0000010010110110","0000001100011001","0000000010011000","1111110111101010","1111101111010100","1111100111110101","1111011111111010","1111011001111001","1111010110001011","1111010000010000","1111000110101010","1110111111010110","1110111110100011","1110111111000000","1110111010101000","1110110101101001","1110111000111010","1111000100010001","1111001110110001","1111010011001010","1111010100011110","1111010111001011","1111011100011101","1111100100101100","1111101111110011","1111111010101001","0000000001101001","0000000110100111","0000001110100100","0000011001010101","0000100001001001","0000100011111001","0000100110110010","0000101110000110","0000110110100000","0000111010001101","0000111000111111","0000110111011110","0000111000111001","0000111100101100","0001000000001111","0001000000101010","0000111100110111","0000110111100110","0000110101001101","0000110101010101","0000110001101100","0000100110010011","0000010111101100","0000001100111111","0000000101111010","1111111100010010","1111101110101110","1111100011011111","1111011111001011","1111011101111101","1111011001101011","1111010010100000","1111001100100010","1111000111101010","1111000000010101","1110111000011101","1110111000000110","1111000001100010","1111001010110111","1111001010000101","1111000011101000","1111000100110000","1111010000100010","1111011011111011","1111011110101001","1111011110011010","1111100011111111","1111101101110101","1111110101011100","1111111100000011","0000000111101110","0000010110110101","0000100001001000","0000100100100101","0000100111101110","0000101110000000","0000110011010001","0000110101010000","0000111000011000","0000111110101101","0001000010010011","0000111111000000","0000111010101111","0000111100100111","0001000000011010","0000111100010010","0000110000011111","0000101000000001","0000101000100010","0000101010000110","0000100010100101","0000010011010101","0000000101101110","1111111110000100","1111111000001100","1111101111111010","1111100110101010","1111011111010100","1111011001001101","1111010010010110","1111001011100011","1111000110111101","1111000100011010","1111000010010010","1111000000100000","1111000000000011","1111000000011101","1111000000110011","1111000010010000","1111000110010101","1111001011101010","1111001111110000","1111010011001011","1111011000001111","1111011110010110","1111100011100111","1111101001110111","1111110100100010","0000000001000000","0000001000100110","0000001011100110","0000010010011011","0000100000000011","0000101011000010","0000101011011001","0000101000001000","0000101101100101","0000111010011000","0001000001010010","0000111101000100","0000110111010101","0000111001010110","0000111111111010","0001000010110001","0001000000011100","0000111100011011","0000110111001010","0000101110010100","0000100010111011","0000011001001101","0000010011000100","0000001101111111","0000000110010101","1111111011000010","1111101110110000","1111100101110101","1111100010000011","1111011111111000","1111011010011100","1111010010000000","1111001011010000","1111001000001000","1111000101110101","1111000010011110","1111000000001100","1111000000100010","1111000001001000","1110111111110110","1110111110101011","1111000001011110","1111001001100011","1111010100101111","1111011110011100","1111100010101000","1111100011001101","1111101000011001","1111110110100110","0000000110000101","0000001100010001","0000001011101101","0000010000100111","0000011101111100","0000101001001101","0000101100010010","0000101110101011","0000110111100000","0001000001101101","0001000101101111","0001000101010000","0001000100010101","0001000000001101","0000110110111100","0000110000001000","0000110010110110","0000111000100111","0000110101110010","0000101010101111","0000100001000101","0000011011001011","0000010010100110","0000000101111001","1111111011110010","1111110111011010","1111110011100000","1111101011101000","1111100010000110","1111011010001000","1111010011100110","1111001110100010","1111001100010010","1111001011000011","1111000110111001","1111000001010011","1111000000110001","1111000110001111","1111001001111100","1111000111010101","1111000101001010","1111001011000111","1111010101010001","1111011010000011","1111011001111011","1111011111000110","1111101101000001","1111111010001000","1111111110000101","1111111110010110","0000000101100011","0000010011010001","0000011101101100","0000100001101001","0000100110101110","0000110001111100","0000111101000100","0001000000100101","0000111111010000","0001000000110110","0001000110000100","0001001000100011","0001000101001010","0000111111010000","0000111010110111","0000111000011001","0000110110011111","0000110011011101","0000101101010110","0000100011111100","0000011010000000","0000010001011011","0000000111111100","1111111011101111","1111110000011010","1111101010011100","1111100111100011","1111100001111001","1111011001010100","1111010011000000","1111010000110101","1111001111100001","1111001101001101","1111001011001011","1111001000110100","1111000011110110","1110111110111101","1111000000010111","1111000111111010","1111001101101001","1111001101101100","1111001110011111","1111010110010011","1111100001000010","1111100111000001","1111101000111101","1111101110010110","1111111001110010","0000000110000101","0000001110100001","0000010100011001","0000011010100110","0000100000111100","0000100101111101","0000101010100110","0000110000110100","0000110111100111","0000111011010100","0000111010011001","0000110111111001","0000110111110101","0000111010010010","0000111011111011","0000111010110011","0000110111111010","0000110011111110","0000101101111111","0000100110001010","0000011110110110","0000011000101001","0000010000111000","0000000110101011","1111111101101001","1111111000000011","1111110010001011","1111101000011101","1111011110100010","1111011001100110","1111010110101111","1111001110111100","1111000011001000","1110111100000011","1110111101010100","1111000001001101","1111000010011100","1111000010011110","1111000011101100","1111000101000110","1111000110110111","1111001011111011","1111010011111000","1111011001110011","1111011100100010","1111100001010001","1111101010110000","1111110100111110","1111111100110011","0000000100101010","0000001101110111","0000010101000100","0000011001111000","0000100001101011","0000101101011010","0000110101101100","0000110111000010","0000111000110110","0001000000011100","0001000110011111","0001000011000011","0000111100000011","0000111100010001","0001000001101011","0001000001011001","0000111001000110","0000110000110001","0000101100011100","0000100111011010","0000011101111000","0000010010011101","0000001000110111","0000000001111111","1111111101101100","1111111010111010","1111110110011101","1111101110011010","1111100101011110","1111011110100001","1111010111011010","1111001101010100","1111000011100111","1111000000000111","1111000010000100","1111000011001011","1111000001010000","1111000000100110","1111000011111101","1111000111111100","1111001001000001","1111001001110100","1111001111101010","1111011010100010","1111100100101110","1111101010101111","1111101111111110","1111111000111101","0000000011100011","0000001010000110","0000001100101111","0000010001101000","0000011010111011","0000100011100010","0000101000100010","0000101110011110","0000111000011010","0001000000110000","0001000010000011","0001000000110110","0001000100011100","0001001010011010","0001001010100110","0001000100100000","0000111111000100","0000111100001101","0000110110000101","0000101001101010","0000011100010100","0000010100011110","0000010001110111","0000001111000110","0000000111101011","1111111011111111","1111110001000010","1111101011001110","1111100111101111","1111011111000110","1111010000101110","1111000110001000","1111000101110000","1111001000111100","1111000110011101","1111000000111010","1111000000111011","1111000101010011","1111000100111101","1110111111011101","1110111110111001","1111000111011000","1111010000101001","1111010100000011","1111010110101101","1111011111000110","1111101001111011","1111110001010100","1111111000000010","0000000100001001","0000010011001110","0000011101011101","0000100010010000","0000101000001100","0000110000101011","0000110101011101","0000110100000100","0000110011000110","0000111000011101","0001000000101000","0001000100100101","0001000010111000","0000111110110111","0000111010101100","0000110111001001","0000110101101111","0000110110010101","0000110100101101","0000101100110111","0000100000001010","0000010011100110","0000001010010100","0000000011111010","1111111101110011","1111110101000100","1111101010000111","1111100010110000","1111100011110011","1111100111011100","1111100001100110","1111010000110010","1111000010010101","1111000000010111","1111000100011010","1111000011011010","1110111110111000","1110111111011111","1111000100101110","1111000110010011","1111000011101001","1111000101010100","1111001110101011","1111011000110000","1111011101110100","1111100001000010","1111100111011111","1111110000101011","1111111001100010","0000000001100111","0000001010011110","0000010100101100","0000011111010110","0000101000011101","0000101110010001","0000110001110001","0000110101111101","0000111010111001","0000111101000010","0000111011111101","0000111100100000","0001000000000111","0001000000000011","0000110111110101","0000101110100100","0000101101011100","0000110001010111","0000101111110000","0000100110101110","0000011101111100","0000011000100111","0000010001010101","0000000101011101","1111111010100101","1111110101011011","1111110010101010","1111101101000111","1111100100111101","1111011101000110","1111010101110000","1111001101110011","1111000110101101","1111000011011111","1111000100010001","1111000101101011","1111000100101010","1111000001111010","1111000000100111","1111000010011100","1111000110010111","1111001011011000","1111010010011000","1111011011010110","1111100011001111","1111101000000011","1111101100100101","1111110011111111","1111111100001101","0000000001101111","0000000110101001","0000001111001010","0000011001010001","0000011111100110","0000100011011101","0000101011000011","0000110101101001","0000111011000111","0000111001100000","0000111000100110","0000111101000001","0001000001000001","0000111111001101","0000111011010111","0000111010011110","0000111001101101","0000110100011100","0000101100110101","0000100111000101","0000100001011110","0000011000011100","0000001110100110","0000001001000101","0000000110100000","0000000000110011","1111110110101010","1111101100100100","1111100100111010","1111011101010101","1111010100010000","1111001100001111","1111001000000010","1111000110110101","1111000101101100","1111000010111111","1110111111110010","1110111110101111","1111000001100010","1111000110010111","1111001001100000","1111001010001101","1111001100001100","1111010010010011","1111011010100000","1111100001111001","1111101001111100","1111110101000010","0000000000000111","0000000101111010","0000001000001101","0000001110110000","0000011011011100","0000100110010000","0000101001010000","0000101010000000","0000110000111001","0000111011111001","0001000001001111","0000111101110010","0000111000101010","0000111000001110","0000111010010011","0000111010000110","0000110111110111","0000110110100011","0000110101001111","0000101111111001","0000100101101101","0000011010111000","0000010011011111","0000001111000101","0000001010011110","0000000100001110","1111111101000101","1111110100110100","1111101001110100","1111011100110001","1111010001110011","1111001011111101","1111001001010111","1111000110011011","1111000010110010","1111000000000100","1110111110001101","1110111100110100","1110111110010111","1111000100101000","1111001011111010","1111001111000000","1111001111001110","1111010010011010","1111011001010001","1111011110110101","1111100010001010","1111101001000110","1111110110100010","0000000100101010","0000001100110011","0000010000001100","0000010101000100","0000011110010100","0000101000111011","0000101111111101","0000110001100111","0000110001011101","0000110101000000","0000111100000000","0000111111011111","0000111100000110","0000111000110010","0000111100110001","0001000010111000","0001000000110000","0000110111001101","0000110000010011","0000101110001110","0000101000011011","0000011011001011","0000001101110001","0000000101101111","1111111111001010","1111110110100101","1111101111101100","1111101100010110","1111100110111111","1111011100111000","1111010100110111","1111010100010011","1111010101010010","1111001111111111","1111000110110111","1111000001010100","1110111111100011","1110111100101100","1110111001010101","1110111010011101","1111000000011010","1111000110011100","1111001010110100","1111010000100100","1111011001011100","1111100011100101","1111101101001011","1111110101101010","1111111100001010","0000000000011101","0000000101001001","0000001100111100","0000010110100000","0000011110010011","0000100100001010","0000101010101011","0000110001110000","0000110101111001","0000110101110010","0000110100111011","0000110110011100","0000111000111100","0000111001100110","0000111001011011","0000111011100000","0000111110100110","0000111101000110","0000110100111010","0000101011110111","0000101000001111","0000100111001000","0000011111111000","0000010000101001","0000000001100101","1111111001011111","1111110101001111","1111101110000011","1111100011110001","1111011011111000","1111011000101110","1111010110111111","1111010010101001","1111001011000010","1111000011000110","1110111111000110","1111000000111010","1111000100110110","1111000101011011","1111000011001011","1111000100001110","1111001010100100","1111010000111000","1111010011101111","1111010111011111","1111011111111110","1111101001010101","1111101111000000","1111110011111000","1111111100001111","0000000101100110","0000001011101101","0000010000111100","0000011001011010","0000100010101010","0000101000100001","0000101101101100","0000110110011100","0000111110110111","0001000000100111","0000111110111000","0001000001011100","0001000110011111","0001000100111101","0000111100010111","0000110101111101","0000110101000011","0000110010001000","0000101000101010","0000011110111010","0000011010100110","0000010111010000","0000001101111110","0000000000011111","1111110101011011","1111101110001011","1111100110111101","1111011110101001","1111011000010011","1111010101001101","1111010010000001","1111001011100010","1111000011010101","1110111101111110","1110111101010010","1110111110101100","1110111111001100","1110111111000010","1111000000000010","1111000010101001","1111000111000101","1111001110110110","1111011001110011","1111100011101100","1111101001000011","1111101100110011","1111110011011101","1111111011000101","1111111110111000","0000000001010100","0000001010000111","0000011001011001","0000100110011011","0000101100111001","0000110010001010","0000111001111001","0000111111000101","0000111101100111","0000111010001000","0000111010000100","0000111011001100","0000111001100011","0000110111010001","0000110111000100","0000110101010011","0000101110001110","0000100110000110","0000100011000010","0000100010101010","0000011101101111","0000010011010101","0000001001000001","0000000001101111","1111111011010001","1111110011011011","1111101010011000","1111100000110000","1111011000001000","1111010011010010","1111010001111011","1111001110111001","1111000111011010","1111000000100100","1111000000010100","1111000100011110","1111000110101100","1111000110011110","1111001000000110","1111001011101100","1111001101011001","1111001101110011","1111010010011000","1111011100000100","1111100101001010","1111101010011111","1111110000001100","1111111001101011","0000000011001010","0000001000100111","0000001110000001","0000011001100101","0000101000001000","0000101111101000","0000101110000011","0000101101011100","0000110101010001","0000111111000000","0001000000011000","0000111011101101","0000111011111001","0001000001110100","0001000001111010","0000110110110011","0000101011001100","0000101010000000","0000101110001011","0000101011100011","0000100001001101","0000010111100010","0000010000100100","0000000110110011","1111111010100001","1111110011011110","1111110011001111","1111110000110011","1111100110001100","1111011001011000","1111010010010110","1111010000000001","1111001100110011","1111000111111110","1111000100000010","1111000000011101","1110111011111000","1110111001100111","1110111101111111","1111000110111000","1111001101100111","1111010000010101","1111010011110110","1111011011011110","1111100011101111","1111100111111110","1111101001111001","1111101111100111","1111111011010000","0000001000000101","0000010000110101","0000010110001011","0000011100010101","0000100100000011","0000101001111000","0000101100100100","0000110000001101","0000111000001001","0001000000111001","0001000011111011","0001000000100100","0000111101000001","0000111101111000","0001000000011000","0000111110111011","0000111000100110","0000110001001001","0000101011011100","0000100110101101","0000100000110111","0000011001001111","0000010000011111","0000000111011011","1111111110011100","1111110101010011","1111101011101000","1111100010011010","1111011100000000","1111011000111110","1111010110000101","1111001111110011","1111000111000011","1111000000010000","1110111101110010","1110111110001111","1110111111110000","1111000001100100","1111000010010000","1111000000110011","1111000000010000","1111000101110111","1111010001010011","1111011011100011","1111100000011111","1111100100101101","1111101101100011","1111111000001111","1111111111000010","0000000011011010","0000001011011010","0000010110111000","0000011111101101","0000100100100010","0000101010110001","0000110011110110","0000111001100001","0000111000101100","0000111000001110","0000111110010000","0001000101000001","0001000010110111","0000111001101011","0000110100111100","0000111000011100","0000111010101101","0000110011100111","0000100111111111","0000100001000000","0000011101111111","0000010110111111","0000001010100011","1111111111111110","1111111011100011","1111111000101100","1111110010010010","1111101010100000","1111100101010011","1111100000011000","1111010110111010","1111001010010110","1111000001011011","1110111110111101","1110111111011100","1110111111100010","1110111111110101","1111000001001011","1111000001111101","1111000001101010","1111000011000000","1111001000100010","1111010001000011","1111011001010111","1111011111100011","1111100011111001","1111101000100110","1111110001001010","1111111110110110","0000001101001101","0000010101110001","0000011000100111","0000011101000111","0000100111101001","0000110010110001","0000110110100011","0000110011110010","0000110010011000","0000110110001101","0000111011011100","0000111110000000","0000111111010111","0001000001111011","0001000011001101","0000111110110101","0000110101110010","0000101110000110","0000101010111110","0000101000101010","0000100010000110","0000010111101101","0000001101101100","0000000101010110","1111111011111110","1111110000011000","1111100101010010","1111011101010000","1111010111111100","1111010100101000","1111010011111111","1111010100100100","1111010001110011","1111001001111110","1111000010000000","1110111111010100","1111000000101001","1111000001100110","1111000010010011","1111000101111111","1111001100001111","1111010001101100","1111010110000110","1111011011100111","1111100001010010","1111100100110111","1111101000110001","1111110001101100","1111111110000101","0000000111111100","0000001110110010","0000010111111000","0000100011011100","0000101010110100","0000101100001010","0000101110110000","0000110111001010","0000111111011010","0001000000110101","0000111110110110","0001000000100010","0001000100111001","0001000101000101","0000111111000101","0000110111011100","0000110010000010","0000101110011101","0000101010100001","0000100100000110","0000011010001001","0000001110111110","0000000111010010","0000000011101001","1111111110000100","1111110001110101","1111100011000010","1111011010000110","1111011001001010","1111011010001001","1111010110010100","1111001101001111","1111000100011011","1111000001011100","1111000011011110","1111000011101101","1110111110010111","1110111001100010","1110111101100011","1111000111110110","1111001101101110","1111001100111110","1111001111111100","1111011100101100","1111101010001100","1111101110000100","1111101101000010","1111110011101110","0000000011010010","0000010000001010","0000010010110010","0000010001000010","0000010100111011","0000100000011001","0000101100100110","0000110010100000","0000110010011101","0000110011100001","0000111010110111","0001000100011110","0001000111100110","0001000010001101","0000111010101000","0000110101101010","0000110001011100","0000101100011101","0000101001101111","0000101001101101","0000100110010000","0000011011110100","0000010000000011","0000001001001001","0000000100000001","1111111011000001","1111110000100010","1111101010100011","1111100111011011","1111100000110001","1111010110101010","1111001110111010","1111001010100010","1111000100111000","1110111101011101","1110111001101111","1110111011111100","1110111111101101","1111000001110101","1111000100100010","1111001001011011","1111001101100101","1111001111010010","1111010010010100","1111011010011011","1111100101000011","1111101101000110","1111110010011100","1111111001011000","0000000011100111","0000001101101101","0000010100010010","0000011000101100","0000011110110110","0000100111101110","0000110000010110","0000110101101010","0000110111110001","0000111000101101","0000111001111010","0000111100001101","0001000000001100","0001000100100101","0001000101101111","0001000001100110","0000111010110011","0000110100110111","0000101110110111","0000100110000011","0000011100001110","0000010101110001","0000010001011010","0000001000110100","1111111011100100","1111110001111011","1111110000101001","1111110000101010","1111101001000010","1111011100001011","1111010011011101","1111010000111001","1111001101110100","1111000110110110","1111000000111001","1111000000010001","1111000001110010","1111000000101100","1110111110100001","1111000000011100","1111000111010010","1111001110101011","1111010011010100","1111010111000001","1111011101011001","1111100110101111","1111101111110101","1111110110100100","1111111100111110","0000000110001110","0000010001100101","0000011010111010","0000100000110000","0000100110101111","0000101111011111","0000110111010100","0000111001001001","0000110111000111","0000111001000000","0001000001010010","0001001001001011","0001001010000010","0001000101101010","0001000001011010","0000111101001001","0000110101001010","0000101010110000","0000100011110111","0000100010000100","0000100000010100","0000011010011101","0000010001001001","0000000101101110","1111111000100010","1111101101001011","1111101000100100","1111100111111101","1111100010000010","1111010100111111","1111001011000100","1111001011000110","1111001101011110","1111001000110000","1111000000110011","1110111110101110","1111000001100000","1111000010100010","1111000011010011","1111001000110010","1111001110100100","1111001101001100","1111001010010111","1111010010011001","1111100011001101","1111101110100100","1111110001010110","1111110110101111","0000000010000001","0000001000100000","0000000111011000","0000001100101100","0000011111110010","0000110001100010","0000110010001001","0000101001110111","0000101100010000","0000111010111001","0001000101011110","0001000010111111","0000111100001011","0000111011100011","0000111111101110","0001000000111011","0000111100010101","0000110101011001","0000101111101111","0000101011001110","0000100100101010","0000011001111000","0000001101000111","0000000011001111","1111111101111000","1111111001011101","1111110010111001","1111101100000111","1111101000001000","1111100101000001","1111011110000011","1111010010111111","1111001001011100","1111000101111111","1111000110100100","1111000101111111","1111000010111110","1111000001000110","1111000011000100","1111000110110111","1111001001000110","1111001001110111","1111001100000100","1111010001011001","1111011001000010","1111100001110111","1111101011000111","1111110011010101","1111111001011001","1111111111000110","0000000111110011","0000010011101010","0000011110001010","0000100011000011","0000100011100100","0000100101000101","0000101011001000","0000110011101011","0000111001100110","0000111010010111","0000111000011011","0000111000001011","0000111011001101","0000111111001110","0001000000101101","0000111101011011","0000110101110010","0000101100110111","0000100101110000","0000011111111001","0000011000011110","0000010000001001","0000001011000101","0000001000101100","0000000001010111","1111110010010011","1111100101001010","1111100010110110","1111100011110111","1111011010010100","1111001000101010","1110111111101101","1111000101001101","1111001011110000","1111001000100010","1111000010001110","1111000010100001","1111000110010111","1111000110110100","1111000110101111","1111001011111100","1111010011011011","1111010111100100","1111011011001010","1111100010110110","1111101010010110","1111101100010001","1111101110011111","1111111001110011","0000001001101000","0000010001110101","0000010010010101","0000010110110100","0000100011010100","0000101110111011","0000110011010000","0000110100100001","0000110111010000","0000111001010100","0000111001000111","0000111001111000","0000111100010010","0000111011001100","0000110100100110","0000101110000100","0000101011111001","0000101010011101","0000100101010010","0000011110011000","0000011001001010","0000010011111010","0000001100000100","0000000100011010","0000000000001111","1111111011101110","1111110000000000","1111011110001111","1111001111110010","1111001010100111","1111001010011010","1111000111110110","1111000010100011","1110111111110100","1111000001001001","1111000001101010","1110111110100110","1110111101000001","1111000010110000","1111001100100111","1111010001110111","1111010000101011","1111010000011010","1111010110110111","1111100001110001","1111101100111000","1111110111111111","0000000011001111","0000001011011000","0000001110110000","0000010001001100","0000010110100111","0000011101101000","0000100011110101","0000101010110010","0000110011110110","0000111011011011","0000111110010000","0000111111101000","0001000011110001","0001000111100000","0001000100101000","0000111100100010","0000110110110110","0000110110101101","0000110111110111","0000110110010111","0000110010010011","0000101011101101","0000100001000101","0000010011110010","0000001000101110","0000000010011011","1111111110000011","1111110111010011","1111101100101001","1111011111011001","1111010011000010","1111001100001101","1111001100000001","1111001100101101","1111000111111011","1111000000000110","1110111101001101","1111000000000001","1111000000010110","1110111011000100","1110111000111100","1111000001001100","1111001101000101","1111010010000100","1111010010110110","1111011010110110","1111101010101010","1111110110010000","1111111000000101","1111111001100010","0000000011001101","0000001111111100","0000010110111010","0000011001111000","0000100000000001","0000101001001110","0000110000001000","0000110100000001","0000110111100100","0000111001101111","0000111001001001","0000111010010110","0001000000111011","0001000110000100","0001000000111110","0000110101111101","0000110001001010","0000110011011110","0000110001110011","0000100111101111","0000011101011100","0000011000000100","0000010001101101","0000000101101110","1111111001010000","1111110001110011","1111101100101110","1111100110010100","1111100000010101","1111011100000101","1111010110011011","1111001110111000","1111001010010101","1111001001100000","1111000101100011","1110111100001010","1110110110000011","1110111010001011","1111000010100011","1111000110000001","1111000101111111","1111001001011000","1111001111110100","1111010011110001","1111010101111110","1111011100110110","1111101001110010","1111110110101010","1111111110100010","0000000011011111","0000001010100010","0000010101010111","0000100001000000","0000101001010110","0000101101011111","0000110000011000","0000110100101001","0000111001000101","0000111011010100","0000111011101110","0000111011011000","0000111001010011","0000110101110110","0000110101010101","0000111001001101","0000111010010000","0000110001110010","0000100101010000","0000011111010011","0000011111011001","0000011011011100","0000010000110111","0000000111110001","0000000011100000","1111111100011110","1111101110010001","1111100000101101","1111011011101110","1111011011011011","1111010111000010","1111001101100111","1111000100101101","1110111111110010","1110111110101111","1111000000101011","1111000011000110","1111000010000101","1110111110001001","1110111101100001","1111000011101011","1111001011110100","1111010000100000","1111010011101000","1111011001101000","1111100001000101","1111100110011111","1111101100110101","1111111010000001","0000001011101101","0000011000000111","0000011011011110","0000011101000011","0000100100000011","0000101110000010","0000110100111011","0000111000111000","0000111101100000","0001000001001010","0000111110011110","0000110110010011","0000110000110011","0000110010110001","0000110111110011","0000111001001100","0000110101111101","0000110001000101","0000101011100110","0000100100101001","0000011100011111","0000010100011001","0000001101000100","0000000111001110","0000000011001011","1111111110100101","1111110101111001","1111101001101101","1111011111000101","1111011000010010","1111010001111111","1111001010000011","1111000011101110","1111000001000110","1110111110100101","1110111010001101","1110111001011010","1111000000011100","1111001001000100","1111001010110110","1111001001000010","1111001101111111","1111011010000010","1111100010001100","1111100001000010","1111011111000001","1111100110001111","1111110101111011","0000000110011001","0000010010111000","0000011010110011","0000011110110011","0000100001001111","0000100110000101","0000101110001100","0000110101110101","0000111010100100","0000111110010110","0001000010000011","0001000001110110","0000111100001000","0000110111010110","0000111010101111","0001000011010010","0001000110100110","0000111111101000","0000110011001101","0000100111111110","0000011111100111","0000011001000000","0000010100000011","0000010000000110","0000001001111111","1111111111000111","1111110001110001","1111100111111010","1111100100110010","1111100100101000","1111100000010001","1111010101001101","1111001000110001","1111000001110101","1111000000101101","1111000000011001","1110111110110100","1110111110110011","1111000001101010","1111000100011000","1111000101010111","1111000111100110","1111001100100001","1111010000100110","1111010010011111","1111010111111011","1111100100101011","1111110001111101","1111110111101000","1111111001110111","0000000011000110","0000010010110011","0000011101111110","0000100001011101","0000100110100111","0000110010001111","0000111011011010","0000111010010101","0000110101101001","0000110111010101","0000111100100110","0000111100000111","0000110110011101","0000110100101110","0000111000111111","0000111011100001","0000110111100111","0000110001001000","0000101011110001","0000100101010100","0000011011011100","0000010000100010","0000000111011111","1111111111100110","1111110111011011","1111101111101011","1111101001010101","1111100011110110","1111011110011111","1111011000010110","1111001111111010","1111000110010000","1111000000101100","1111000010011010","1111000110010000","1111000101011001","1111000001111010","1111000010100100","1111000101111101","1111000100111100","1111000001100110","1111000111000110","1111010110111110","1111100011110111","1111100101011111","1111100101110110","1111110001000011","0000000010001110","0000001100000101","0000001101100101","0000010001000101","0000011010011110","0000100010111001","0000100101111000","0000101000011111","0000110000101000","0000111100010010","0001000100011100","0001000101001011","0001000001000001","0000111101110001","0000111110100011","0001000000110010","0001000000001010","0000111100000101","0000110110100110","0000101111110000","0000100111000011","0000011111010111","0000011010101110","0000010100000111","0000000110001111","1111110111000011","1111110001100101","1111110100010001","1111110010000111","1111100111011001","1111011110100100","1111011100011101","1111010111100110","1111001010101001","1111000000100010","1111000011000001","1111001010001000","1111001001110011","1111000100110111","1111000100110011","1111001000001100","1111000111111010","1111000110100101","1111001100000010","1111010110010011","1111011101001000","1111100000100101","1111100111010010","1111110001011111","1111111010010101","0000000010011111","0000001101100001","0000010111101110","0000011011010000","0000011100100110","0000100100111101","0000110010010011","0000111001110111","0000111001011010","0000111001001010","0000111100111010","0001000000010100","0001000001101101","0001000011100011","0001000010110001","0000111001011010","0000101100001010","0000100111000010","0000101010010101","0000101001000000","0000011101110001","0000010010111101","0000001111101100","0000001011101110","1111111110110000","1111101111001100","1111100111011001","1111100110001000","1111100011110110","1111011110111101","1111011001011011","1111010001111000","1111001000011101","1111000011010111","1111000101100101","1111000111011000","1111000001111100","1110111011111100","1110111111101110","1111001010001111","1111001111100110","1111001101101110","1111001110011010","1111010111100110","1111100011111001","1111101100010110","1111110001000001","1111110101111101","1111111101101011","0000001000010110","0000010100000000","0000011101000111","0000100010000100","0000100101011001","0000101001101011","0000101101100000","0000101111100001","0000110010110010","0000111010000011","0001000001011011","0001000010101011","0000111110101100","0000111100001111","0000111101111111","0000111111000100","0000111010010111","0000110001000111","0000101000101011","0000100100000001","0000100000011011","0000011000111011","0000001101000100","0000000010101111","1111111110001111","1111111010101001","1111110000010100","1111100001101110","1111011001001110","1111011000111111","1111010111000011","1111001101010001","1111000011000011","1111000000110010","1111000010111111","1111000010000101","1110111111010000","1110111111111111","1111000011001100","1111000100101111","1111000110110100","1111001101100110","1111010101111000","1111011001101111","1111011011001101","1111100000100111","1111101001011011","1111110000111010","1111111000101100","0000000101101010","0000010100101111","0000011101111100","0000100001100011","0000100111000010","0000101111100011","0000110100110111","0000110101111101","0000111000100011","0000111101001111","0000111101111111","0000111010100111","0000111010100101","0000111111001011","0000111111111110","0000111001011101","0000110011010001","0000110010010100","0000110000001011","0000100111010111","0000011101011110","0000011000101001","0000010100010111","0000001010010010","1111111110000101","1111110110101000","1111110001101011","1111101000110110","1111011110000000","1111010111110001","1111010101011101","1111010000101111","1111001001010100","1111000100110010","1111000011101011","1111000000011101","1110111001110000","1110110101010110","1110110111101001","1110111110111000","1111000111111101","1111010001101110","1111011010011010","1111011111011011","1111100001101010","1111100101100000","1111101100111011","1111110101011000","1111111100111100","0000000101010000","0000001111111001","0000011010111101","0000100011010010","0000101000001011","0000101011110000","0000110000011110","0000110110101000","0000111011011011","0000111100010011","0000111011100010","0000111110100111","0001000101100011","0001001000001000","0001000000011111","0000110100111101","0000110000010110","0000110010011100","0000110000011111","0000100101011010","0000011000011010","0000010000101011","0000001010111010","0000000001010000","1111110110011111","1111110000111100","1111101110011000","1111100110100101","1111011001001011","1111001111101101","1111001111110011","1111010011010001","1111010001111101","1111001100101000","1111001000000101","1111000011101000","1110111100010001","1110110110001000","1110111000101101","1111000010011110","1111001001011000","1111001001111000","1111001100001111","1111010110111110","1111100100001101","1111101011011111","1111101111000100","1111110110111001","0000000010111011","0000001100100001","0000010011000010","0000011100100101","0000101001110001","0000110010100010","0000110010101111","0000110001011000","0000110110100001","0000111111101110","0001000100001100","0001000000110111","0000111011010100","0000111010000111","0000111101100011","0001000000001101","0000111100110010","0000110011101101","0000101010010001","0000100011110100","0000011101110111","0000010101000110","0000001011101011","0000000101110100","0000000010000111","1111111011100110","1111110010001100","1111101010100011","1111100101101100","1111011111100110","1111010111001011","1111010000001111","1111001100000010","1111000111011001","1111000010010010","1111000001011011","1111000101010011","1111000111000100","1111000011100011","1111000001011001","1111000110100001","1111001110000111","1111010000011111","1111001111100001","1111010011100101","1111011110110011","1111101011011011","1111110100111101");

begin
   process(RESET,SA_CLK)
   begin
      if RESET = '1' then
         datax <= (others=>'0');
         datad <= (others=>'0');
      elsif rising_edge(SA_CLK) then
         sdatax <= sdatax(1 to len-1) & sdatax(0);
         sdatad <= sdatad(1 to len-1) & sdatad(0);
         datax(ex_wx-1 downto ex_wx-wx) <= sdatax(0);
         datax(ex-1 downto 0) <= (others=>'0');
         datad(ex_wx-1 downto ex_wx-wx) <= sdatad(0);
         datad(ex-1 downto 0) <= (others=>'0');
      end if;
   end process;
end behavioural;
--===========================================================--
--=================== Clock divider =========================--
--===========================================================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;

entity Clock_divider is
   port (
      CLOCK_50 : in  std_logic;
      FCLK     : out std_logic; -- Folding frequency
      XCLK     : out std_logic; -- Main/external clock 12.5MHz
      SA_CLK   : out std_logic; -- 48.828 kHz
      BCLK     : out std_logic; -- XCLK/4 = 3.125 MHz
      SCLK     : out std_logic);-- SPI clock, choose 6.25 MHz
                                -- for timing requirements
end entity Clock_divider;

architecture Behavioural of Clock_divider is

   signal count_SA : integer range 0 to 512 := 0;
   signal count_B  : integer range 0 to 8 := 0;
   signal count_F  : integer range 0 to 5 := 0;
   signal count_X  : integer range 0 to 2 := 0;
   signal count_S  : integer range 0 to 4 := 0;
   signal sSA_CLK  : std_logic := '0';
   signal sBCLK    : std_logic := '0';
   signal sSCLK    : std_logic := '0';
   signal sXCLK    : std_logic := '0';
   signal sFCLK    : std_logic := '0';

begin
   SA_CLK   <= sSA_CLK;
   BCLK     <= sBCLK;
   SCLK     <= sSCLK;
   XCLK     <= sXCLK;
   FCLK     <= sFCLK;
   process(CLOCK_50)
   begin
      if rising_edge(CLOCK_50) then
         count_F <= count_F + 1;
         count_B <= count_B + 1;
         count_X <= count_X + 1;
         count_S <= count_S + 1;
         count_SA <= count_SA + 1;
         if count_B = 7 then -- CLOCK_50/16 = 3.125 MHz
            count_B <= 0;
            sBCLK <= not(sBCLK);
         end if;
         --Clock divider 12.5MHz---------------------
         if count_X = 1 then -- CLOCK_50/4 = 12.5 MHz
            count_X <= 0;
            sXCLK <= not(sXCLK);
         end if;
         --Clock divider 6.25 MHz--------------------
         if count_S = 3 then -- CLOCK_50/8 = 6.25 MHz
            count_S <= 0;
            sSCLK <= not(sSCLK);
         end if;
         --Clock divider 48.828 kHz------------------
         if count_SA = 511 then -- CLOCK_50/1024 = 48.828 kHz
            sSA_CLK <= not(sSA_CLK);
            count_SA <= 0;
         end if;
         if count_F = 512/fl - 1 then
            sFCLK <= not(sFCLK);
            count_F <= 0;
         end if;
      end if;
   end process;
end Behavioural;

--===========================================================--
--=================== Audio interface =======================--
--===========================================================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;

entity Audio_Interface is
   port(
      CLOCK_IN  : in  std_logic;  -- Sampling clock for DAC
      CLOCK_OUT : in  std_logic;  -- Sampling clock for ADC
      BCLK      : in  std_logic;  -- Bit clock
      DIN       : out std_logic;  -- Data bit in to AIC23
      DOUT      : in  std_logic;  -- Data bit out from AIC23
      -- For processing --
      ADC_L     : out byte_data;  -- Data register from AIC23, channel left
      ADC_R     : out byte_data;  -- Data register from AIC23, channel right
      DAC_L     : in  byte_data;  -- Data register to AIC23, channel left
      DAC_R     : in  byte_data); -- Data register to AIC23, channel right
end Audio_Interface;

architecture Behavioural of Audio_Interface is

signal get_L : byte_data:=(others=>'0');
signal get_R : byte_data:=(others=>'0');
signal count_inL  : natural range 0 to 100 := 0;
signal count_inR  : natural range 0 to 100 := 0;
signal count_outL : natural range 0 to 100 := 0;
signal count_outR : natural range 0 to 100 := 0;

begin
   --Counting for sampling the audio data
   process(BCLK)
   begin
      if falling_edge(BCLK) then
         count_outL <= count_outL + 1;
         count_outR <= count_outR + 1;
         count_inL <= count_inL + 1;
         count_inR <= count_inR + 1;
      -- output channel -----
         case CLOCK_OUT is
            when '0'=>count_outR <= 0;
                        ADC_R <= get_R;
            when '1'=>count_outL <= 0;
                        ADC_L <= get_L;
            when others=>null;
         end case;
      -- input channel ------
         case CLOCK_IN is
            when '0'=>count_inR <= 0;
            when '1'=>count_inL <= 0;
            when others=>null;
         end case;
      -----------------------
      end if;
   end process;
   --Input the audio signals
   process(BCLK)
   begin
      if rising_edge(BCLK) then
         if (count_outL>0) and (count_outL<wx+2) then
            get_L <= get_L(wx-2 downto 0) & DOUT;
         end if;
         if (count_outR>0) and (count_outR<wx+2) then
            get_R <= get_R(wx-2 downto 0) & DOUT;
         end if;
      end if;
   end process;
   --Output the audio signals
   DIN <= DAC_L(wx - count_inL) when (count_inL>0) and (count_inL<wx+1) else
          DAC_R(wx - count_inR) when (count_inR>0) and (count_inR<wx+1) else
          '0';
end Behavioural;
--===========================================================--
--=================== Audio controller ======================--
--===========================================================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;

entity Audio_Controller is
   port(
      CLOCK_50   : in  std_logic;
      SCLK       : in  std_logic;  -- SPI clock
      AIC_SPI_CS : out std_logic;  -- SPI CS, ack for new command
      AD_SDIO    : out std_logic;  -- SPI data
      I2C_SCLK   : out std_logic;  -- I2C clock
      I2C_SDAT   : out std_logic); -- I2C data
end entity Audio_Controller;

architecture Behavioural of Audio_Controller is
   --====SPI controller====--
   signal position_SPI : natural range 0 to 18 := 0;
   signal list_CMD     : natural range 0 to 12 := 0;

   subtype CMD_type is std_logic_vector(0 to 15);
   signal COMMAND : CMD_type;
   --Left/right line inputs : 0dB, normal
   constant LLI_vol     : CMD_type := "0000000"&"01"&"00"&"10111";
   constant RLI_vol     : CMD_type := "0000001"&"01"&"00"&"10111";
   --Left/right headphone outputs : 0dB, no zero-cross detect
   constant LHI_vol     : CMD_type := "0000010"&"00"&"1111001";
   constant RHI_vol     : CMD_type := "0000011"&"00"&"1111001";
   --Analogue path: No sidetone, disable mic, ADC : line inputs
   constant ana_path    : CMD_type := "0000100"&"000"&"010"&"100";
   --Digital path: 48kHz
   constant dig_path    : CMD_type := "0000101"&"00000"&"0110"; -- ??? should enable HPF?
   --Power down: no power down
   constant PWR_down    : CMD_type := "0000110"&"000000001";
   --Master/16bit/I2S
   constant dif_format  : CMD_type := "0000111"&"001000010";
   --MCLK/48/256fs/Normal
   constant sam_rate    : CMD_type := "0001000"&"000000000";
   --Activate
   constant dif_activ   : CMD_type := "0001001"&"000000001";
   --Write 000000000
   constant rset_reg    : CMD_type := "0001111"&"000000000";
   --====I2C controller====--
   signal sI2C_SCLK: std_logic := '1';
   signal sI2C_SDAT: std_logic := '1';
   signal count_I  : integer range 0 to 132 := 0;
   signal I2C_pos  : natural range 0 to 30 := 0;
   signal I2C_COMMAND : CMD_type;
   signal I2C_list_CMD: natural range 0 to 12 := 0;
   type I2C_Mstate is (idle,start_I2C,stop_I2C,trans_I2C);
   signal state_I2C,nstate_I2C : I2C_Mstate := idle;
   constant ini_RW : std_logic_vector(0 to 7) := "00110100";
begin
--================SPI controller=====================--
--Command pulse process--------------------------------
AD_SDIO <= COMMAND(position_SPI) when position_SPI < 16
           else '1';
--SPI Creating commands positions process----
   SPI_pos: process(SCLK)
   begin
      if falling_edge(SCLK) then
         position_SPI <= position_SPI + 1;
         if list_CMD < 12 then
            AIC_SPI_CS <= '0';
         else
            AIC_SPI_CS <= '1';
         end if;
         if position_SPI = 15 then
            if list_CMD < 12 then
               list_CMD <= list_CMD + 1;
               AIC_SPI_CS <= '1';
            end if;
         elsif position_SPI = 16 then
            position_SPI <= 0;
         end if;
      end if;
   end process;
--SPI Audio mode process--------------------
   SPI_mode: process(SCLK)
   begin
      if rising_edge(SCLK) then
         case list_CMD is
            when 0=>COMMAND <= rset_reg;
            when 1=>COMMAND <= rset_reg;
            when 2=>COMMAND <= LLI_vol;
            when 3=>COMMAND <= RLI_vol;
            when 4=>COMMAND <= LHI_vol;
            when 5=>COMMAND <= RHI_vol;
            when 6=>COMMAND <= ana_path;
            when 7=>COMMAND <= dig_path;
            when 8=>COMMAND <= PWR_down;
            when 9=>COMMAND <= dif_format;
            when 10=>COMMAND <= sam_rate;
            when 11=>COMMAND <= dif_activ;
            when others=>COMMAND <= (others=> '1'); 
         end case;
      end if;
   end process;
--================I2C controller=====================--
   I2C_SCLK <= sI2C_SCLK;
   I2C_SDAT <= ini_RW(I2C_pos-1) when (I2C_pos>0) and (I2C_pos<9) else
               I2C_COMMAND(I2C_pos-10) when (I2C_pos>9) and (I2C_pos<18) else
               I2C_COMMAND(I2C_pos-11) when (I2C_pos>18) and (I2C_pos<27) else
               sI2C_SDAT;
   with I2C_list_CMD select
   I2C_COMMAND <= rset_reg   when 0,
                  LLI_vol    when 1,
                  RLI_vol    when 2,
                  LHI_vol    when 3,
                  RHI_vol    when 4,
                  ana_path   when 5,
                  dig_path   when 6,
                  PWR_down   when 7,
                  dif_format when 8,
                  sam_rate   when 9,
                  dif_activ  when 10,
                  (others=> '1') when others;
--State machine--
   FSM_I2C: process(nstate_I2C)
   begin
      state_I2C <= nstate_I2C;
   end process;
--I2S Creating commands positions process----
   I2C_position_creation: process(CLOCK_50)
   begin
      if rising_edge(CLOCK_50) then
         if I2C_list_CMD < 11 then
            count_I <= count_I + 1;
         end if;
         if (state_I2C /= idle) and (state_I2C /= stop_I2C) then
            if count_I = 30 then
               I2C_pos <= I2C_pos + 1;
            elsif count_I = 65 then -- CLOCK_50/132 = 378.79 kHz
               sI2C_SCLK <= '1';
            elsif count_I = 131 then
               sI2C_SCLK <= '0';
               count_I <= 0;
            end if;
         end if;
         -- I2C interface ----------------------------------
         case state_I2C is
            -- Prepare for starting ------------------
            when idle=>
               if count_I < 80 then
                  sI2C_SCLK <= '1';
                  sI2C_SDAT <= '1';
               else
                  nstate_I2C <= start_I2C;
               end if;
            -- Create starting condition -------------
            when start_I2C=>
               sI2C_SDAT <= '0';
               if count_I = 65 then
                  nstate_I2C <= trans_I2C;
               end if;
            -- Position for sending command ----------
            when trans_I2C=>
               if I2C_pos = 28 then
                  I2C_pos <= 0;
                  nstate_I2C <= stop_I2C;
                  count_I <= 0;
               end if;
            -- Create stopping condition -------------
            when stop_I2C=>
               if (count_I<20) then
                  sI2C_SCLK <= '0';
               elsif (count_I<70) then
                  sI2C_SCLK <= '1';
                  sI2C_SDAT <= '0';
               else
                  if I2C_list_CMD < 11 then
                     I2C_list_CMD <= I2C_list_CMD + 1;
                     nstate_I2C <= idle;
                  end if;
               end if;
         end case;         
      end if;
   end process;
--I2C Sending commands ---------------------
end Behavioural;

--===========================================================--
--=================== FIR filter direct form I ==============--
--===========================================================--

--=================== DIRECT FORM I PE ======================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;
--library lpm;
use work.LPM_COMPONENTS.all;

entity PE_DI is
   port(
      RESET  : in    std_logic;
      SA_CLK : in    std_logic;
      XIN    : in    byte_exdata; -- Input to PE
      HIN    : in    byte_exdata; -- Coefficient to PE
      YIN    : in    byte_exproduct; -- Output to PE
      EIN    : in    byte_exdata; -- Error to be multiplied to XIN

      XOUT   : inout byte_exdata; -- Input from PE
      YOUT   : out   byte_exproduct; -- Output from PE
      EXOUT  : out   byte_exproduct);-- EIN*XIN
end entity PE_DI;

architecture DI_FIR_behav of PE_DI is

signal pr: byte_exproduct := (others => '0');

begin
   -- Flip flop 1 --
   FF_1: LPM_FF
      generic map(
         LPM_WIDTH=> ex_wx)
      port map (
         DATA    => XIN,
         CLOCK   => SA_CLK,
         ACLR    => RESET,
         ENABLE  => '1',
         Q       => XOUT);
   -- Multiplier 1 --------
   MULT_1: LPM_MULT
      GENERIC MAP (
         LPM_WIDTHA=> ex_wx, LPM_WIDTHB=> ex_wx, 
         LPM_REPRESENTATION=>"SIGNED", 
         LPM_WIDTHP=> ex_wp, 
         LPM_WIDTHS=> ex_wp)  
      PORT MAP (
         DATAA => XOUT,
         DATAB => HIN,
         RESULT=> pr);
   -- Adder 1 -------------
   ADD_1: LPM_ADD_SUB
      GENERIC MAP (
         LPM_WIDTH => ex_wp,
         LPM_REPRESENTATION=>"SIGNED",
         LPM_DIRECTION=>"ADD")
      PORT MAP (
         DATAA => pr,
         DATAB => YIN,
         RESULT=> YOUT);
   -- Calculate EXOUT = e*x*mu --
   CAL: LPM_MULT   -- Multiply xemu(i) = emu * x(i)
      GENERIC MAP(
         LPM_WIDTHA=> ex_wx, LPM_WIDTHB=> ex_wx, 
         LPM_REPRESENTATION=>"SIGNED", 
         LPM_WIDTHP=> ex_wp, 
         LPM_WIDTHS=> ex_wp)
      PORT MAP(
         DATAA => XIN,
         DATAB => EIN, 
         RESULT=> EXOUT);
end DI_FIR_behav;

--======== NORMAL FIR filter direct form I ==================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;

entity FIR_DI is
   port(
      RESET  : in  std_logic;
      SA_CLK : in  std_logic;
      XIN    : in  byte_exdata; -- Filter input
      EIN    : in  byte_exdata; -- Error in
      YOUT   : out byte_exproduct; -- Filter output

      HIN    : in  array_exdata; -- Filter coefficient
      EXOUT  : out array_exproduct);-- e*x
end FIR_DI;

architecture Behavioural of FIR_DI is

signal sYOUT  : byte_exproduct :=(others=>'0');
signal datay  : array_exproduct:=(others=>(others=>'0'));
signal datax  : array_exdata:=(others=>(others=>'0'));
begin
----FIR filter--------------------------------------------
   -- First PE ---------------
   PE_first: PE_DI
   port map(
      RESET   => RESET,
      SA_CLK  => SA_CLK,
      XIN     => XIN,         -- First Xin
      HIN     => HIN(fl-1),   -- First Hin
      YIN     => datay(fl-1), -- First Yin
      EIN     => EIN,         -- First Ein

      Xout    => datax(fl-2), -- Second Xin
      YOUT    => datay(fl-2), -- Second Yin
      EXOUT   => EXOUT(fl-1));-- Second Ein
   -- Create middle PEs -------
   PE_loop: for i in (fl-2) downto 1 generate
   PE_middle: PE_DI
   port map(
      RESET  => RESET,
      SA_CLK => SA_CLK,
      XIN    => datax(i), 
      HIN    => HIN(i),   
      YIN    => datay(i),
      EIN    => EIN,

      XOUT   => datax(i-1),
      YOUT   => datay(i-1),
      EXOUT  => EXOUT(i));
   end generate;
   -- Last PE ----------------
   PE_last: PE_DI
   port map(
      RESET  => RESET,
      SA_CLK => SA_CLK,
      XIN    => datax(0),
      HIN    => HIN(0),
      YIN    => datay(0),
      EIN    => EIN,
      
      YOUT   => sYOUT,
      EXOUT  => EXOUT(0));
----------------------------------------------------------
   YOUT <= sYOUT;
end Behavioural;

--============ FOLDING FIR direct form I ====================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;
--library lpm;
use work.LPM_COMPONENTS.all;

entity FIR_DI_FOLDING is
   port(
      RESET   : in  std_logic;
      CLOCK_F : in  std_logic;
      XIN     : in  byte_exdata; -- Filter input
      EIN     : in  byte_exdata; -- Error in
      YOUT    : out byte_exproduct; -- Filter output

      HIN     : in  array_exdata; -- Filter coefficient
      EXOUT   : out array_exproduct);-- e*x
end FIR_DI_FOLDING;

architecture Behavioural of FIR_DI_FOLDING is

signal sxin   : array_exdata    := (others=>(others=>'0'));
signal cntCR  : natural range 0 to 1024 := 0;
signal DR     : array_DR        := (others=>(others=>'0'));
signal pr     : byte_exproduct  := (others=>'0');
signal addr   : byte_exproduct  := (others=>'0');
signal sYOUT  : byte_exproduct  := (others=>'0');
signal outmux : byte_exproduct  := (others=>'0');
signal outff  : byte_exproduct  := (others=>'0');
signal shin   : byte_exdata     := (others=>'0');

signal EXOUT_2d : array_exproduct := (others=>(others=>'0'));
signal sEXOUT : byte_exproduct  := (others=>'0');

begin
   --Coefficients shifted out--
   --EXOUT <= sEXOUT;
   shin <= Hin(fl-1-cntCR);
   YOUT <= sYOUT;
   --Create coefficients register position--
   process(RESET,CLOCK_F)
   begin
      if RESET = '1' then
         cntCR <= 0;
      elsif rising_edge(CLOCK_F) then
         cntCR <= cntCR + 1;
         --SR block--
         DR <= DR(fl-1 downto 0) & DR(fl);
         if cntCR = fl-1 then
            cntCR <= 0;
         --CR block--
            sxin <= XIN & sxin(fl-1 downto 1);
            DR(fl) <= sxin(fl-1);
            sYOUT <= addr;
         end if;
      end if;
   end process;
   --Flip flop--
   FF_1: LPM_FF
      generic map(
         LPM_WIDTH=> ex_wp)
      port map (
         DATA    => outmux,
         CLOCK   => CLOCK_F,
         ACLR    => RESET,
         ENABLE  => '1',
         Q       => outff);
   --Multiplier block--
   Multiplier: lpm_mult --multr = h*x
   GENERIC MAP(
      LPM_WIDTHA=> ex_wx, LPM_WIDTHB=> ex_wx,
      LPM_REPRESENTATION=>"SIGNED",
      LPM_WIDTHP=> ex_wp,
      LPM_WIDTHS=> ex_wp)
   PORT MAP(
      dataa => DR(fl),
      datab => shin,
      result=> pr);
   --Adder block--
   Adder: LPM_ADD_SUB --addr = pr + outmux
   GENERIC MAP(
      LPM_WIDTH => ex_wp,
      LPM_REPRESENTATION=>"SIGNED",
      LPM_DIRECTION=>"ADD")
   PORT MAP(
      DATAA => pr,
      DATAB => outff,
      RESULT=> addr);
   --MUX-------
   outmux <= addr when cntCR < fl-1 else
             (others=>'0');
   -- Calculate EXOUT = e*x*mu--
   CAL_EXMU: for i in fl - 1 downto 0 generate
   MULT_1: LPM_MULT   --Multiply xemu(i) = emu * x(i)
      GENERIC MAP(
         LPM_WIDTHA=> ex_wx, LPM_WIDTHB=> ex_wx,
         LPM_REPRESENTATION=>"SIGNED",
         LPM_WIDTHP=> ex_wp,
         LPM_WIDTHS=> ex_wp)
      PORT MAP(
         DATAA => sxin(i),
         DATAB => EIN,
         RESULT=> EXOUT(i));
   end generate;
end Behavioural;

--============ LMS ADF FOLDING DI ===========================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;
--library lpm;
use work.LPM_COMPONENTS.all;

entity FIR_DI_FOLDING_LMS is
   port(
      RESET   : in  std_logic;
      CLOCK_F : in  std_logic;
      SA_CLK  : in  std_logic;
      XIN     : in  byte_exdata; -- Primary signal
      DIN     : in  byte_exdata; -- Desired signal
      EOUT    : out byte_exdata; -- error out
      YOUT    : out byte_exdata);-- filter output
end FIR_DI_FOLDING_LMS;

architecture Behavioural of FIR_DI_FOLDING_LMS is

--Adaptive FIR filter
   --Array of coefficients
   signal hin_2d  : array_exdata:=(others=>(others=>'0')); 
   signal exmu    : array_exproduct:=(others=>(others=>'0'));
   
   signal sxdin   : byte_exproduct:=(others=>'0'); --Size extension
   signal sxyout  : byte_exproduct:=(others=>'0');
   signal seout   : byte_exproduct:=(others=>'0');
   signal syout   : byte_exproduct:=(others=>'0');
   signal emu     : byte_exdata:=(others=>'0');
   
begin
--Interface-------------------------------------------------
   eout <= seout(ex_wx downto 1);
   yout <= sxyout(ex_wx-1 downto 0);
--Initialization --
   --Signed extension to product length---------------------
   sxdin(ex_wx-1 downto 0) <= din;
   sxdin(ex_wp-1 downto ex_wx) <= (others=>din(din'high)); --Signed extension
   --Rearrange the output to after being multiplied---------
   sxyout(ex_wx-1 downto 0) <= syout(ex_wp-1-fx downto ex_wx-fx); --Extract the data value
   sxyout(ex_wp-1 downto ex_wx) <= (others=>syout(syout'high)); --Signed extension
   --Calculate the error and emu ---------------------------
   seout <= sxdin - sxyout; -- could be round up to 1 bit
   emu <= seout(ex_wx-1+4 downto 4); -- Divided by 2^4
   --Update the coefficients--------------------------------
   process(SA_CLK)
   begin
      if rising_edge(SA_CLK) then
         for i in fl-1 downto 0 loop
            hin_2d(i) <= hin_2d(i) + exmu(i)(ex_wp-1-fx+4 downto ex_wx-fx+4); --Divided by 2^4
         end loop;
      end if;
   end process;
   --FIR filter---------------------------------------------
   FIR_DI_FOLDING_block: FIR_DI_FOLDING
   port map(
      RESET    => RESET,
      CLOCK_F  => CLOCK_F,
      XIN      => xin,
      HIN      => hin_2d,
      EIN      => emu,

      YOUT     => syout,
      EXOUT    => exmu);
end Behavioural;

--============== LMS ADF filter direct form I ===============--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;
--library lpm;
use work.LPM_COMPONENTS.all;

entity LMS_ADF_DI is
  port (
      RESET   : in  std_logic;      
      SA_CLK  : in  std_logic;
      XIN     : in  byte_exdata; -- Primary signal
      DIN     : in  byte_exdata; -- Desired signal
      EOUT    : out byte_exdata; -- error out
      YOUT    : out byte_exdata);-- filter output
end LMS_ADF_DI;

architecture Behavioural of LMS_ADF_DI is
--Adaptive FIR filter
   --Array of coefficients
   signal hin_2d  : array_exdata:=(others=>(others=>'0')); 
   signal exmu    : array_exproduct:=(others=>(others=>'0'));
   
   signal sxdin   : byte_exproduct:=(others=>'0'); --Size extension
   signal sxyout  : byte_exproduct:=(others=>'0');
   signal seout   : byte_exproduct:=(others=>'0');
   signal syout   : byte_exproduct:=(others=>'0');
   signal emu     : byte_exdata:=(others=>'0');
   
begin
--Interface-------------------------------------------------
   eout <= seout(ex_wx-1 downto 0);
   yout <= sxyout(ex_wx-1 downto 0);
--Initialization --
   --Signed extension to product length---------------------
   sxdin(ex_wx-1 downto 0) <= din;
   sxdin(ex_wp-1 downto ex_wx) <= (others=>din(din'high)); --Signed extension
   --Rearrange the output to after being multiplied---------
   sxyout(ex_wx-1 downto 0) <= syout(ex_wp-1-fx downto ex_wx-fx); --Extract the data value
   sxyout(ex_wp-1 downto ex_wx) <= (others=>syout(syout'high)); --Signed extension
   --Calculate the error and emu ---------------------------
   seout <= sxdin - sxyout;
   emu <= seout(ex_wx-1+4 downto 4); -- Divided by 2^4
   --Update the coefficients--------------------------------
   process(SA_CLK)
   begin
      if rising_edge(SA_CLK) then
         for i in fl-1 downto 0 loop
            hin_2d(i) <= hin_2d(i) + exmu(i)(ex_wp-1-fx+4 downto ex_wx-fx+4); --Divided by 2^4
         end loop;
      end if;
   end process;
   --FIR filter---------------------------------------------
   FIR_DI_block: FIR_DI
   port map(
      SA_CLK => SA_CLK,
      RESET  => RESET,
      XIN    => XIN,
      HIN    => HIN_2d,
      EIN    => emu,

      YOUT   => sYOUT,
      EXOUT  => exmu);
end Behavioural;
--===========================================================--
--============== FIR filter direct form II ==================--
--===========================================================--

--=================== DIRECT FORM II PE =====================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;
--library lpm;
use work.LPM_COMPONENTS.all;

entity PE_DII is
   port (
      RESET  : in    std_logic;
      SA_CLK : in    std_logic;
      XIN    : in    byte_exdata; -- Input to PE
      HIN    : in    byte_exdata; -- Coefficient to PE
      YIN    : in    byte_exproduct; -- Output to PE
      EIN    : in    byte_exdata; -- Error to be multiplied to XIN
      
      XOUT   : inout byte_exdata; -- Input from PE
      YOUT   : out   byte_exproduct; -- Output from PE
      EXOUT  : out   byte_exproduct);-- EIN*XIN
end entity PE_DII;

architecture DII_FIR_behav of PE_DII is

signal pr: byte_exproduct := (others => '0');
signal su: byte_exproduct := (others => '0');

begin
   XOUT <= XIN;
   -- Multiplier 1 --------
   MULT_1: LPM_MULT
      GENERIC MAP (
         LPM_WIDTHA=> ex_wx, LPM_WIDTHB=> ex_wx, 
         LPM_REPRESENTATION=>"SIGNED", 
         LPM_WIDTHP=> ex_wp, 
         LPM_WIDTHS=> ex_wp)  
      PORT MAP(
         DATAA => XIN,
         DATAB => HIN,
         RESULT=> pr);
   -- Adder 1 -------------
   ADD_1: LPM_ADD_SUB
      GENERIC MAP (
         LPM_WIDTH => ex_wp,
         LPM_REPRESENTATION=>"SIGNED",
         LPM_DIRECTION=>"ADD")
      PORT MAP(
        DATAA => pr,
        DATAB => YIN,
        RESULT=>su);
   -- Flip flop 1 --
   FF_1: LPM_FF
      GENERIC MAP (
         LPM_WIDTH=> ex_wp)
      PORT MAP(
         DATA    =>su,
         CLOCK   => SA_CLK,
         ACLR    => RESET,
         ENABLE  => '1',
         Q       => YOUT);
   -- Calculate EXOUT = e*x*mu--
   CAL: LPM_MULT   --Multiply xemu(i) = emu * x(i)
      GENERIC MAP(
         LPM_WIDTHA=> ex_wx, LPM_WIDTHB=> ex_wx, 
         LPM_REPRESENTATION=>"SIGNED", 
         LPM_WIDTHP=> ex_wp, 
         LPM_WIDTHS=> ex_wp)
      PORT MAP(
         DATAA => XIN,
         DATAB => EIN, 
         RESULT=> EXOUT);
end DII_FIR_behav;

--======= NORMAL FIR filter direct form II ==================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;

entity FIR_DII is
   port(
      RESET  : in  std_logic;
      SA_CLK : in  std_logic;
      XIN    : in  byte_exdata; -- Filter input
      EIN    : in  byte_exdata; -- Error in
      YOUT   : out byte_exproduct; -- Filter output

      HIN    : in  array_exdata; -- Filter coefficient
      EXOUT  : out array_exproduct);-- e*x
end FIR_DII;

architecture Behavioural of FIR_DII is

signal sYOUT : byte_exproduct:=(others=>'0');
signal datay : array_exproduct:=(others=>(others=>'0'));
signal datax : array_exdata:=(others=>(others=>'0'));

begin
----FIR filter--------------------------------------------
   -- First PE ---------------
   PE_first: PE_DII
   port map(
      RESET => RESET,
      SA_CLK=> SA_CLK,
      XIN   => XIN,         -- First Xin
      HIN   => HIN(0),      -- First Hin
      YIN   => datay(fl-1), -- First Yin
      EIN   => EIN,         -- First Ein

      XOUT  => datax(fl-2), -- Second Xin
      YOUT  => datay(fl-2), -- Second Yin
      EXOUT => EXOUT(fl-1));-- Second Ein
   -- Create middle PEs -------
   PE_loop: for i in (fl-2) downto 1 generate
   PE_middle: PE_DII
   port map(
      RESET  => RESET,
      SA_CLK => SA_CLK,
      XIN    => datax(i),
      HIN    => HIN(fl-1-i),
      YIN    => datay(i),
      EIN    => EIN,

      XOUT   => datax(i-1),
      YOUT   => datay(i-1),
      EXOUT  => EXOUT(i));
   end generate;
   -- Last PE ----------------
   PE_last: PE_DII
   port map(
      RESET  => RESET,
      SA_CLK => SA_CLK,
      XIN    => datax(0),
      HIN    => HIN(fl-1),
      YIN    => datay(0),
      EIN    => EIN,
      
      YOUT   => sYOUT,
      EXOUT  => EXOUT(0));
----------------------------------------------------------
   YOUT <= sYOUT;
end Behavioural;

--============ FOLDING FIR direct form II ===================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;
--library lpm;
use work.LPM_COMPONENTS.all;

entity FIR_DII_FOLDING is
   port(
      RESET   : in  std_logic;
      CLOCK_F : in  std_logic;
      XIN     : in  byte_exdata; -- Filter input
      EIN     : in  byte_exdata; -- Error in
      YOUT    : out byte_exproduct; -- Filter output

      HIN     : in  array_exdata; -- Filter coefficient
      EXOUT   : out array_exproduct);-- e*x
end FIR_DII_FOLDING;

architecture Behavioural of FIR_DII_FOLDING is

signal sxin   : array_exdata    := (others=>(others=>'0'));
signal cntCR  : natural range 0 to fl - 1 := fl - 1;
signal SR     : array_SR := (others=>(others=>'0'));
signal pr     : byte_exproduct  := (others=>'0');
signal addr   : byte_exproduct  := (others=>'0');
signal shin   : byte_exdata     := (others=>'0');
signal outmux : byte_exproduct  := (others=>'0');

begin
   --Coefficients shifted out--
   shin <= Hin(fl-1-cntCR);
   --Create coefficients register position--
   process(RESET,CLOCK_F)
   begin
      if RESET = '1' then
         cntCR <= fl - 1;
      elsif rising_edge(CLOCK_F) then
         --SR block--
         SR <= addr & SR(fl downto 1);
         --CR block--
         if cntCR = 0 then
            cntCR <= fl - 1;
            sxin <= XIN & sxin(fl-1 downto 1);
         else
            cntCR <= cntCR - 1;
         end if;
         --Output--
         if cntCR = fl-1 then
            YOUT <= SR(fl);
         end if;
      end if;
   end process;
   --Multiplier block--
   Multiplier: lpm_mult --multr = h*x
   GENERIC MAP(
      LPM_WIDTHA=> ex_wx, LPM_WIDTHB=> ex_wx,
      LPM_REPRESENTATION=>"SIGNED",
      LPM_WIDTHP=> ex_wp,
      LPM_WIDTHS=> ex_wp)
   PORT MAP(
      dataa => sxin(fl-1),
      datab => shin,
      result=> pr);
   --Adder block--
   Adder: LPM_ADD_SUB --addr = pr + outmux
   GENERIC MAP(
      LPM_WIDTH => ex_wp,
      LPM_REPRESENTATION=>"SIGNED",
      LPM_DIRECTION=>"ADD")
   PORT MAP(
      DATAA => pr,
      DATAB => outmux,
      RESULT=> addr);
   --MUX-------
   outmux <= (others=>'0') when cntCR = fl-1 else
             SR(0);
   -- Calculate EXOUT = e*x*mu--
   CAL_EXMU: for i in fl - 1 downto 0 generate
   MULT_1: LPM_MULT   --Multiply xemu(i) = emu * x(i)
      GENERIC MAP(
         LPM_WIDTHA=> ex_wx, LPM_WIDTHB=> ex_wx,
         LPM_REPRESENTATION=>"SIGNED",
         LPM_WIDTHP=> ex_wp,
         LPM_WIDTHS=> ex_wp)
      PORT MAP(
         DATAA => sxin(i),
         DATAB => EIN,
         RESULT=> EXOUT(i));
   end generate;
end Behavioural;

--============== LMS ADF filter direct form II ==============--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;
--library lpm;
use work.LPM_COMPONENTS.all;

entity LMS_ADF_DII is
  port (
      RESET   : in  std_logic;      
      SA_CLK  : in  std_logic;
      XIN     : in  byte_exdata; -- Primary signal
      DIN     : in  byte_exdata; -- Desired signal
      EOUT    : out byte_exdata; -- error out
      YOUT    : out byte_exdata);-- filter output
end LMS_ADF_DII;

architecture Behavioural of LMS_ADF_DII is
--Adaptive FIR filter
   --Array of coefficients
   signal hin_2d : array_exdata:=(others=>(others=>'0'));
   signal exmu   : array_exproduct:=(others=>(others=>'0'));
   
   signal sxdin  : byte_exproduct:=(others=>'0'); --Size extension
   signal sxyout : byte_exproduct:=(others=>'0');
   signal seout  : byte_exproduct:=(others=>'0');
   signal syout  : byte_exproduct:=(others=>'0');
   signal emu    : byte_exdata:=(others=>'0');
   
begin
--Interface-------------------------------------------------
   eout <= seout(ex_wx-1 downto 0);
   yout <= sxyout(ex_wx-1 downto 0);
--Initialization --
   --Signed extension to product length---------------------
   sxdin(ex_wx-1 downto 0) <= din;
   sxdin(ex_wp-1 downto ex_wx) <= (others=>din(din'high)); --Signed extension
   --Rearrange the output to after being multiplied---------
   sxyout(ex_wx-1 downto 0) <= syout(ex_wp-1-fx downto ex_wx-fx); --Extract the data value
   sxyout(ex_wp-1 downto ex_wx) <= (others=>syout(syout'high)); --Signed extension
   --Calculate the error and emu ---------------------------
   seout <= sxdin - sxyout;
   emu <= seout(ex_wx-1+4 downto 4); -- Divided by 2^4
   --Update the coefficients--------------------------------
   process(SA_CLK)
   begin
      if rising_edge(SA_CLK) then
         for i in fl-1 downto 0 loop
            hin_2d(i) <= hin_2d(i) + exmu(i)(ex_wp-1-fx+4 downto ex_wx-fx+4); --Divided by 2^4
         end loop;
      end if;
   end process;
   --FIR filter---------------------------------------------
   FIR_DII_block: FIR_DII
   port map(
      SA_CLK => SA_CLK,
      RESET  => RESET,
      XIN    => XIN,
      HIN    => HIN_2d,
      EIN    => emu,
      YOUT   => sYOUT,
      EXOUT  => exmu);
end Behavioural;

--============ LMS ADF FOLDING DII ==========================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;
--library lpm;
use work.LPM_COMPONENTS.all;

entity FIR_DII_FOLDING_LMS is
   port(
      RESET   : in  std_logic;      
      CLOCK_F : in  std_logic;
      SA_CLK  : in  std_logic;
      XIN     : in  byte_exdata; -- Primary signal
      DIN     : in  byte_exdata; -- Desired signal
      EOUT    : out byte_exdata; -- error out
      YOUT    : out byte_exdata);-- filter output
end FIR_DII_FOLDING_LMS;

architecture Behavioural of FIR_DII_FOLDING_LMS is

--Adaptive FIR filter
   --Array of coefficients
   signal hin_2d  : array_exdata:=(others=>(others=>'0')); 
   signal exmu    : array_exproduct:=(others=>(others=>'0'));
   
   signal sxdin   : byte_exproduct:=(others=>'0'); --Size extension
   signal sxyout  : byte_exproduct:=(others=>'0');
   signal seout   : byte_exproduct:=(others=>'0');
   signal syout   : byte_exproduct:=(others=>'0');
   signal emu     : byte_exdata:=(others=>'0');

begin
--Interface-------------------------------------------------
   eout <= seout(ex_wx downto 1);
   yout <= sxyout(ex_wx-1 downto 0);
--Initialization --
   --Signed extension to product length---------------------
   sxdin(ex_wx-1 downto 0) <= din;
   sxdin(ex_wp-1 downto ex_wx) <= (others=>din(din'high)); --Signed extension
   --Rearrange the output to after being multiplied---------
   sxyout(ex_wx-1 downto 0) <= syout(ex_wp-1-fx downto ex_wx-fx); --Extract the data value
   sxyout(ex_wp-1 downto ex_wx) <= (others=>syout(syout'high)); --Signed extension
   --Calculate the error and emu ---------------------------
   seout <= sxdin - sxyout;
   emu <= seout(ex_wx-1+4 downto 4); -- Divided by 2^5
   --Update the coefficients--------------------------------
   process(SA_CLK)
   begin
      if rising_edge(SA_CLK) then
         for i in fl-1 downto 0 loop
            hin_2d(i) <= hin_2d(i) + exmu(i)(ex_wp-1-fx+4 downto ex_wx-fx+4); --Divided by 2^5
         end loop;
      end if;
   end process;
   --FIR filter---------------------------------------------
   FIR_DII_FOLDING_block: FIR_DII_FOLDING
   port map(
      RESET    => RESET,
      CLOCK_F  => CLOCK_F,
      XIN      => xin,
      HIN      => hin_2d,
      EIN      => emu,

      YOUT     => syout,
      EXOUT    => exmu);
end Behavioural;

--===========================================================--
--============ FOLDING FIR direct form I 50MHZ ==============--
--===========================================================--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.my_pack.all;
--library lpm;
use work.LPM_COMPONENTS.all;

entity FIR_DI_FOLDING_50MHz is
   port(
      RESET    : in  std_logic;
      CLOCK_50 : in  std_logic;
      XIN      : in  byte_exdata; -- Filter input
      EIN      : in  byte_exdata; -- Error in
      YOUT     : out byte_exproduct; -- Filter output

      HIN      : in  array_exdata; -- Filter coefficient
      EXOUT    : out array_exproduct);-- e*x
end FIR_DI_FOLDING_50MHz;

architecture Behavioural of FIR_DI_FOLDING_50MHz is

signal sxin   : array_exdata    := (others=>(others=>'0'));
signal cntCR  : natural range 0 to 1024 := 0;
signal posCR  : natural range 0 to fl := 0;
signal DR     : array_DR        := (others=>(others=>'0'));
signal pr     : byte_exproduct  := (others=>'0');
signal addr   : byte_exproduct  := (others=>'0');
signal outmux : byte_exproduct  := (others=>'0');
signal outff  : byte_exproduct  := (others=>'0');
signal shin   : byte_exdata     := (others=>'0');

begin
   --Coefficients shifted out--
   shin <= Hin(fl-1-posCR);
   posCR <= cntCR when (cntCR < fl) else
            0;
   --Create coefficients register position--
   process(RESET,CLOCK_50)
   begin
      if RESET = '1' then
         cntCR <= 0;
      elsif rising_edge(CLOCK_50) then
         cntCR <= cntCR + 1;
         if cntCR < fl then
            if cntCR = fl-1 then
               YOUT <= addr;
            end if;
         --DR block--
            DR <= DR(fl-1 downto 0) & DR(fl);
         elsif cntCR = 1023 then
            sxin <= XIN & sxin(fl-1 downto 1);
            DR(fl) <= sxin(fl-1);
            cntCR <= 0;
         else
            DR(fl) <= (others => '0');
         end if;
      end if;
   end process;
   --Flip flop--
   FF_1: LPM_FF
      generic map(
         LPM_WIDTH=> ex_wp)
      port map (
         DATA    => outmux,
         CLOCK   => CLOCK_50,
         ACLR    => RESET,
         ENABLE  => '1',
         Q       => outff);
   --Multiplier block--
   Multiplier: lpm_mult --multr = h*x
   GENERIC MAP(
      LPM_WIDTHA=> ex_wx, LPM_WIDTHB=> ex_wx,
      LPM_REPRESENTATION=>"SIGNED",
      LPM_WIDTHP=> ex_wp,
      LPM_WIDTHS=> ex_wp)
   PORT MAP(
      dataa => DR(fl),
      datab => shin,
      result=> pr);
   --Adder block--
   Adder: LPM_ADD_SUB --addr = pr + outmux
   GENERIC MAP(
      LPM_WIDTH => ex_wp,
      LPM_REPRESENTATION=>"SIGNED",
      LPM_DIRECTION=>"ADD")
   PORT MAP(
      DATAA => pr,
      DATAB => outff,
      RESULT=> addr);
   --MUX-------
   outmux <= addr when cntCR < fl-1 else
             (others=>'0');
   -- Calculate EXOUT = e*x*mu--
   CAL_EXMU: for i in fl - 1 downto 0 generate
   MULT_1: LPM_MULT   --Multiply xemu(i) = emu * x(i)
      GENERIC MAP(
         LPM_WIDTHA=> ex_wx, LPM_WIDTHB=> ex_wx,
         LPM_REPRESENTATION=>"SIGNED",
         LPM_WIDTHP=> ex_wp,
         LPM_WIDTHS=> ex_wp)
      PORT MAP(
         DATAA => sxin(i),
         DATAB => EIN,
         RESULT=> EXOUT(i));
   end generate;
end Behavioural;